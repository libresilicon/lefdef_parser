VERSION 5.7 ;
# DEMO4 CHIP - 1280 ARRAY

#&alias &&area = (73600,74400) (238240,236400) &endalias
#&alias &&core = (85080,85500) (226760,224700) &endalias
#&alias &&m2stripes = sroute stripe net vss net vdd layer m2
#    width
#    320 count 2 pattern 87900 4200 218100
#    area &&area core &&core &endalias
#&alias &&m3stripes = sroute stripe net vss net vdd layer m3
#    width
#    600 count 2 pattern 89840 6720 217520 area
#    &&area core &&core &endalias
#&alias &&powerfollowpins = sroute follow net vss net vdd layer
#    m1 width 560
#    area &&area core &&core &endalias
#&alias &&powerrepair = sroute repair net vss net vdd area
#    &&area core &&core &endalias
# PLACEMENT SITE SECTION

LAYER POLYS
  TYPE MASTERSLICE ;
END POLYS

LAYER PW
  TYPE MASTERSLICE ;
END PW

LAYER NW
  TYPE MASTERSLICE ;
END NW

LAYER PD
  TYPE MASTERSLICE ;
END PD

LAYER ND
  TYPE MASTERSLICE ;
END ND

LAYER CUT01
  TYPE CUT ;
END CUT01

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 5.6 ;
  WIDTH2.6 ;
  SPACING 1.5 ;
END M1

LAYER CUT12
  TYPE CUT ;
END CUT12

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 6.0 ;
  WIDTH 3.2 ;
  SPACING 1.6 ;
END M2

LAYER CUT23
  TYPE CUT ;
END CUT23

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 5.6 ;
  WIDTH 3.6;
  SPACING 1.6 ;
END M3

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA C2PW DEFAULT
  LAYER PW ;
  RECT -2.0 -2.0 2.0 2.0 ;
  LAYER CUT01 ;
  RECT -0.6 -0.6 0.6 0.6 ;
  LAYER M1 ;
  RECT -2.0 -2.0 2.0 2.0 ;
END C2PW

VIA C2NW DEFAULT
 LAYER NW ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT01 ;
 RECT -0.6 -0.6 0.6 0.6 ;
 LAYER M1 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END C2NW

VIA C2PD DEFAULT
 LAYER PD ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT01 ;
 RECT -0.6 -0.6 0.6 0.6 ;
 LAYER M1 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END C2PD

VIA C2ND DEFAULT
 LAYER ND ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT01 ;
 RECT -0.6 -0.6 0.6 0.6 ;
 LAYER M1 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END C2ND

VIA C2POLY DEFAULT
 LAYER POLYS ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT01 ;
 RECT -0.6 -0.6 0.6 0.6 ;
 LAYER M1 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END C2POLY

VIA VIA12 DEFAULT
 LAYER M1 ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT12 ;
 RECT -0.7 -0.7 0.7 0.7 ;
 LAYER M2 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END VIA12

VIA VIA23 DEFAULT LAYER M3 ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT23 ;
 RECT -0.8 -0.8 0.8 0.8 ;
 LAYER M2 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END VIA23

SPACING SAMENET
  CUT01 CUT12 4.0 ;
  SAMENET CUT12 CUT23 4.0 ;
END SPACING

VIA VIACENTER12 LAYER M1 ;
 RECT -4.6 -2.2 4.6 2.2 ;
 LAYER CUT12 ;
 RECT -3.1 -0.8 -1.9 0.8 ;
 RECT 1.9 -0.8 3.1 0.8 ;
 LAYER M2 ;
 RECT -4.4 -2.0 4.4 2.0 ;
END VIACENTER12

VIA VIATOP12
 LAYER M1 ;
 RECT -2.2 -2.2 2.2 8.2 ;
 LAYER CUT12 ;
 RECT -0.8 5.2 0.8 6.8 ;
 LAYER M2 ;
 RECT -2.2 -2.2 2.2 8.2 ;
END VIATOP12

VIA VIABOTTOM12 LAYER M1 ;
 RECT -2.2 -8.2 2.2 2.2 ;
 LAYER CUT12 ;
 RECT -0.8 -6.8 0.8 -5.2 ;
 LAYER M2 ;
 RECT -2.2 -8.2 2.2 2.2 ;
END VIABOTTOM12

VIA VIALEFT12 LAYER M1 ;
 RECT -7.8 -2.2 2.2 2.2 ;
 LAYER CUT12 ;
 RECT -6.4 -0.8 -4.8 0.8 ;
 LAYER M2 ;
 RECT -7.8 -2.2 2.2 2.2 ;
END VIALEFT12

VIA VIARIGHT12
 LAYER M1 ;
 RECT -2.2 -2.2 7.8 2.2 ;
 LAYER CUT12 ;
 RECT 4.8 -0.8 6.4 0.8 ;
 LAYER M2 ;
 RECT -2.2 -2.2 7.8 2.2 ;
END VIARIGHT12

VIA VIABIGPOWER12 LAYER M1 ;
 RECT -21.0 -21.0 21.0 21.0 ;
 LAYER CUT12 ;
 RECT -2.4 -0.8 2.4 0.8 ;
 RECT -19.0 -19.0 -14.2 -17.4 ;
 RECT -19.0 17.4 -14.2 19.0;
 RECT 14.2 -19.0 19.0 -17.4 ;
 RECT 14.2 17.4 19.0 19.0 ;
 RECT -19.0 -0.8 -14.2 0.8 ;
 RECT -2.4 -19.0 2.4 -17.4 ;
 RECT 14.2 -0.8 19 0.8 ;
 RECT -2.4 17.4 2.4 19.0 ;
 LAYER M2 ;
 RECT -21.0 -21.0 21.0 21.0 ;
END VIABIGPOWER12

VIARULE VIALIST12
 LAYER M1 ;
 DIRECTION VERTICAL ;
 WIDTH 9.0 TO 9.6;
 LAYER M2 ;
 DIRECTION HORIZONTAL ;
 WIDTH 3.0 TO 3.0 ;
 VIA VIACENTER12 ;
 VIA VIATOP12 ;
 VIA VIABOTTOM12 ;
 VIA VIALEFT12 ;
 VIA VIARIGHT12 ;
END VIALIST12

VIARULE VIAGEN12 GENERATE LAYER M1 ;
 ENCLOSURE 0.01 0.05 ;
 LAYER M2 ;
 ENCLOSURE 0.01 0.05 ;
 LAYER CUT12 ;
 RECT -0.06 -0.06 0.06 0.06 ;
 SPACING 0.14 BY 0.14 ;
 END VIAGEN12 VIA VIACENTER23 LAYER M3 ;
 RECT -2.2 -2.2 2.2 2.2 ;
 LAYER CUT23 ;
 RECT -0.8 -0.8 0.8 0.8 ;
 LAYER M2 ;
 RECT -2.0 -2.0 2.0 2.0 ;
 END VIACENTER23 VIA VIATOP23 LAYER M3 ;
 RECT -2.2 -2.2 2.2 8.2 ;
 LAYER CUT23 ;
 RECT -0.8 5.2 0.8 6.8 ;
 LAYER M2 ;
 RECT -2.2 -2.2 2.2 8.2 ;
END VIATOP23

VIA VIABOTTOM23 LAYER M3 ;
 RECT -2.2 -8.2 2.2 2.2 ;
 LAYER CUT23 ;
 RECT -0.8 -6.8 0.8 -5.2 ;
 LAYER M2 ;
 RECT -2.2 -8.2 2.2 2.2 ;
END VIABOTTOM23

VIA VIALEFT23
 LAYER M3 ;
 RECT -7.8 -2.2 2.2 2.2 ;
 LAYER CUT23 ;
 RECT -6.4 -0.8 -4.8 0.8 ;
 LAYER M2 ;
 RECT -7.8 -2.2 2.2 2.2 ;
END VIALEFT23

VIA VIARIGHT23
 LAYER M3 ;
 RECT -2.2 -2.2 7.8 2.2 ;
 LAYER CUT23 ;
 RECT 4.8 -0.8 6.4 0.8 ;
 LAYER M2 ;
 RECT -2.2 -2.2 7.8 2.2 ;
END VIARIGHT23

VIARULE VIALIST23
 LAYER M3 ;
 DIRECTION VERTICAL ;
 WIDTH 3.6 TO 3.6 ;
 LAYER M2 ;
 DIRECTION HORIZONTAL ;
 WIDTH 3.0 TO 3.0 ;
 VIA VIACENTER23 ;
 VIA VIATOP23 ;
 VIA VIABOTTOM23 ;
 VIA VIALEFT23 ;
 VIA VIARIGHT23 ;
END VIALIST23

VIARULE VIAGEN23 GENERATE
 LAYER M2 ;
 ENCLOSURE 0.01 0.05 ;
 LAYER M3 ;
 ENCLOSURE 0.01 0.05 ;
 LAYER CUT23 ;
 RECT -0.06 -0.06 0.06 0.06 ;
 SPACING 0.14 BY 0.14 ;
END VIAGEN23

#MOVED SIDE BLOCK HERE AS SPECIFIED BY POSITION IN LEFMANUAL
SITE CORE1 SIZE 67.2 BY 6 ; # GCD of all Y sizes of Macros
END CORE1

SITE IOX
  SIZE 37.8 BY 444 ; # 151.2 / 4 = 37.8 , 4 sites per pad
END IOX

SITE IOY
  SIZE 436.8 BY 30 ; # 150 / 5 = 30 , 5 sites per pad
END IOY

SITE SQUAREBLOCK
  SIZE 268.8 BY 252 ;
END SQUAREBLOCK

SITE I2BLOCK
  SIZE 672 BY 504 ;
END I2BLOCK

SITE LBLOCK
  SIZE 201.6 BY 168 ;
END LBLOCK

SITE CORNER
  SIZE 436.8 BY 444 ;
END CORNER

MACRO CORNER
 CLASS ENDCAP BOTTOMLEFT ;
 SIZE 436.8 BY 444 ;
 SYMMETRY X Y ;
 SITE CORNER ;
 PIN VDD SHAPE RING ;
   DIRECTION INOUT ;
   PORT LAYER M2 ;
     WIDTH 20 ;
     PATH 426.8 200 200 200 200 434 ;
   END
 END VDD
 PIN VSS
  SHAPE RING ;
  DIRECTION INOUT ;
  PORT
    LAYER M2 ;
    WIDTH 20 ;
    PATH 100 434 100 100 ;
    LAYER M1;
    WIDTH 20 ;
    PATH 100 100 426.8 100 ;
  END
  END VSS
END CORNER

MACRO IN1X
 class pad ;
 FOREIGN IN1X ;
 SIZE 151.2 BY 444 ;
 SYMMETRY X ;
 SITE IOX ;
 PIN Z DIRECTION OUTPUT ;
   PORT
   LAYER M1 ;
      PATH 61.6 444 72.8 444 ;
   END
 END Z
PIN PO
   DIRECTION OUTPUT ;
   PORT
     LAYER M1 ;
     PATH 78.4 444 84.0 444 ;
   END
  END PO
  PIN A
   DIRECTION INPUT ;
   PORT
      LAYER M1 ;
      PATH 95.2 444 100.8 444 ;
   END
   END A
  PIN PI
   DIRECTION INPUT ;
   PORT
   LAYER M1 ;
   PATH 106.4 444 112 444 ;
  END
 END PI
 PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      WIDTH 20 ;
      PATH 10 200 141.2 200 ;
    END
 END VDD
 PIN VSS
 DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT
   LAYER M1 ;
   WIDTH 20 ;
   PATH 10 100 141.2 100 ;
 END
END VSS
END IN1X

MACRO IN1Y EEQ IN1X ;
 FOREIGN IN1Y ;
 class pad ;
 SIZE 436.8 BY 150 ;
 SYMMETRY Y ;
 SITE IOY ;
 PIN Z DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      PATH 0 69 0 75 ;
    END
 END Z
 PIN PO
    DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      PATH 0 81 0 87 ;
    END
 END PO
 PIN A DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 51 0 57 ;
 END
END A PIN PI DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 39 0 45 ;
 END
END PI PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 236.8 10 236.8 140 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 336.8 10 336.8 140 ;
 END
END VSS
END IN1Y

MACRO FILLER FOREIGN FILLER ;
 SIZE 67.2 BY 6 ;
 SYMMETRY X Y;
 SITE CORE1 ;
 PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M1 ;
 RECT 45.8 0 55 6 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M1 ;
 RECT 12.2 0 21.4 6 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 4.5 ;
 END
END FILLER MACRO INV FOREIGN INVS ;
 SIZE 67.2 BY 24 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 30.8 9 42 9 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 15 ;
 END
END A PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 13.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 13.4 ;
 END

END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 16.5 ;
 END
END INV MACRO BUF FOREIGN BUFS ;
 SIZE 67.2 BY 126 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 39 42 39 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 30.8 33 ;
 END
END A PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 10.0 56.0 10.0 56.0 115.8 50.4 115.8 50.4 121.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 10.0 11.2 10.0 11.2 115.8 16.8 115.8 16.8 121.4 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 124.5 ;
 END
END BUF

MACRO BIDIR1X FOREIGN BIDIR1X ;
 class pad ;
 SIZE 151.2 BY 444 ;
 SYMMETRY X ;
 SITE IOX ;
 PIN IO DIRECTION INOUT ;
 PORT LAYER M1 ;
 PATH 61.6 444 67.2 444 ;
 END
END IO PIN ZI DIRECTION OUTPUT ;
 PORT LAYER M1 ;
 PATH 78.4 444 84.0 444 ;
 END
END ZI PIN PO DIRECTION OUTPUT ;
 PORT LAYER M1 ;
 PATH 95.2 444 100.8 444 ;
 END
END PO PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 106.4 444 112.0 444 ;
 END
END A PIN EN DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 134.4 444 140.0 444 ;
 END
END EN PIN TN DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 28.0 444 33.6 444 ;
 END
END TN PIN PI DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 44.8 444 50.4 444 ;
 END
END PI PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 10 200 141.2 200 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
PORT LAYER M1 ;
 WIDTH 20 ;
 PATH 10 100 141.2 100 ;
 END
END VSS
END BIDIR1X

MACRO BIDIR1Y EEQ BIDIR1X ;
 class pad ;
 FOREIGN BIDIR1Y ;
 SIZE 436.8 BY 150 ;
 SYMMETRY Y ;
 SITE IOY ;
 PIN IO DIRECTION INOUT ;
 PORT LAYER M2 ;
 PATH 0 69 0 75 ;
 END
END IO PIN ZI DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 0 93 0 99 ;
 END
END ZI PIN PO DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 0 81 0 87 ;
 END
END PO PIN A DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 15 0 21 ;
 END
END A PIN EN DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 27 0 33 ;
 END
END EN PIN TN DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 39 0 45 ;
 END
END TN PIN PI DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 51 0 57 ;
 END
END PI PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 236.8 10 236.8 140 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 336.8 10 336.8 140 ;
 END
END VSS
END BIDIR1Y

MACRO OR2
 FOREIGN OR2S ;
 SIZE 67.2 BY 42 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 39 42 39 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 15 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 3 ;
 END
END B PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 10.0 ;
 PATH 50.4 27.4 50.4 37.4 ;
 VIA 50.4 3 C2PW ;
 VIA 50.4 21 C2PW ;
 VIA 50.4 33 C2PW ;
 VIA 50.4 39 C2PW ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 10.0 ;
 PATH 16.8 27.4 16.8 37.4 ;
 VIA 16.8 3 C2NW ;
 VIA 16.8 15 C2NW ;
 VIA 16.8 21 C2NW ;
 VIA 16.8 33 C2NW ;
 VIA 16.8 39 C2NW ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 40.5 ;
 END
END OR2

MACRO AND2 FOREIGN AND2S ;
 SIZE 67.2 BY 84 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 39 42 39 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 42 15 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 42 3 ;
 END
END B PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 79.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 79.4 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 82.5 ;
 END
END AND2

MACRO DFF3
 FOREIGN DFF3S ;
 SIZE 67.2 BY 210 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Q DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 19.6 99 47.6 99 ;
 END
END Q PIN QN DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 123 42 123 ;
 END
END QN PIN D DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 30.8 51 ;
 END
END D PIN G DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 3 ;
 END
END G PIN CD DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 36.4 75 ;
 END
END CD PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 205.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 205.4 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 208.5 ;
 PATH 8.4 3 8.4 123 ;
 PATH 58.8 3 58.8 123 ;
 PATH 64.4 3 64.4 123;
 END
END DFF3

MACRO NOR2
 FOREIGN NOR2S ;
 SIZE 67.2 BY 42 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M1 ;
 PATH 42 33 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 15 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 36.4 9 ;
 END
END B PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 37.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 37.4 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 40.5 ;
 END
END NOR2

MACRO AND2J
 EEQ AND2 ;
 FOREIGN AND2SJ ;
 SIZE 67.2 BY 48 ;
 SYMMETRY X Y ;
 ORIGIN 0 6 ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 33 42 33 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 42 15 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 42 3 ;
 END
END B PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 -1.4 50.4 37.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 -1.4 16.8 37.4 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 34.5 ;
 END
END AND2J

MACRO SQUAREBLOCK FOREIGN SQUAREBLOCKS ;
 CLASS RING ;
SIZE 268.8 BY 252 ;
 SITE SQUAREBLOCK ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 22.8 21 246.0 21 ;
 END
END Z PIN A DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 64.4 33 137.2 33 ;
 PATH 137.2 33 137.2 69 ;
 PATH 137.2 69 204.4 69 ;
 END
END A PIN B DIRECTION INPUT ;
PORT LAYER M2 ;
 PATH 22.8 129 246.0 129 ;
 END
END B PIN C DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 70 165 70 153 ;
 PATH 70 153 126 153 ;
 END
END C PIN D DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 22.8 75 64.4 75 ;
 END
END D PIN E DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 22.8 87 64.4 87 ;
 END
END E PIN F DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 22.8 99 64.4 99 ;
 END
END F PIN G DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 22.8 111 64.4 111 ;
 END
END G PIN VDD DIRECTION INOUT ;
 SHAPE RING ;
 PORT LAYER M1 ;
 WIDTH 3.6 ;
 PATH 4.0 3.5 4.0 248 ;
 PATH 264.8 100 264.8 248 ;
 PATH 150 3.5 150 100 ;
 LAYER M2 ;
 WIDTH 3.6 ;
 PATH 4.0 3.5 150 3.5 ;
 PATH 150 100 264.8 100 ;
 PATH 4.0 248 264.8 248 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE RING ;
 PORT LAYER M1 ;
 WIDTH 3.6 ;
 PATH 10 10 10 150 ;
 PATH 100 150 100 200 ;
 PATH 50 200 50 242 ;
 PATH 258.8 10 258.8 242 ;
 LAYER M2 ;
 WIDTH 3.6 ;
 PATH 10 150 100 150 ;
 PATH 100 200 50 200 ;
 PATH 10 10 258.8 10 ;
 PATH 50 242 258.8 242 ;
 END
END VSS OBS LAYER M1 ;
 RECT 13.8 14.0 255.0 237.2 ;
 END
END SQUAREBLOCK

MACRO I2BLOCK FOREIGN I2BLOCKS ;
 CLASS RING ;
 SIZE 672 BY 504 ;
 SITE I2BLOCK ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 22.8 21 649.2 21 ;
 END
END Z PIN A DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 22.8 63 154.0 63 ;
 PATH 154.0 63 154.0 129;
 PATH 154.0 129 447.6 129 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 137.2 423 447.6 423 ;
 END
END B PIN C DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 204.4 165 271.6 165 ;
 END
END C PIN D DIRECTION INPUT ;
PORT LAYER M2 ;
 PATH 204.4 171 271.6 171 ;
 END
END D PIN E DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 204.4 213 204.4 213 ;
 END
END E PIN F DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 406 249 406 273 ;
 END
END F PIN G DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 338.8 249 338.8 273 ;
 END
END G PIN H DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 372.4 357 372.4 381 ;
 END
END H PIN VDD DIRECTION INOUT ;
 SHAPE RING ;
 PORT LAYER M1 ;
 WIDTH 3.6 ;
 PATH 668 3.5 668 80.5 ;
 PATH 467 80.5 467 465.5 ;
 PATH 668 465.5 668 500.5 ;
 PATH 4 500.5 4 465.5 ;
 PATH 138 465.5 138 80.5 ;
 PATH 4 80.5 4 3.5 ;
 LAYER M2 ;
 WIDTH 3.6 ;
 PATH 4 3.5 668 3.5;
 PATH 668 80.5 467 80.5 ;
 PATH 467 465.5 668 465.5 ;
 PATH 668 500.5 4 500.5 ;
 PATH 4 465.5 138 465.5 ;
 PATH 138 80.5 4 80.5 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE RING ;
 PORT LAYER M1 ;
 WIDTH 3.6 ;
 PATH 662 10 662 74 ;
 PATH 461 74 461 472 ;
 PATH 662 472 662 494 ;
 PATH 10 494 10 472;
 PATH 144 472 144 74 ;
 PATH 10 74 10 10 ;
LAYER M2 ;
 WIDTH 3.6 ;
 PATH 10 10 662 10 ;
 PATH 662 74 461 74 ;
 PATH 461 472 662 472 ;
 PATH 662 494 10 494 ;
 PATH 10 472 144 472 ;
 PATH 144 74 10 74 ;
 END
END VSS OBS LAYER M1 ;
 RECT 14 14 658 70 ;
 RECT 14 476 658 490 ;
 RECT 148 14 457 490 ;
 # rectilinear shape description LAYER OVERLAP ;
 RECT 0 0 672 84 ;
 RECT 134.4 84 470.4 462 ;
 RECT 0 462 672 504 ;
 END
END I2BLOCK

MACRO LBLOCK
 FOREIGN LBLOCKS ;
 CLASS RING ;
 SIZE 201.6 BY 168 ;
 SITE LBLOCK ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 2.8 15 198.8 15 ;
 END
END Z PIN A DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 2.8 81 137.2 81 ;
 PATH 137.2 81 137.2 69 ;
 PATH 137.2 69 198.8 69 ;
 END
END A
PIN B DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 2.8 165 64.4 165 ;
 END
END B PIN C DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 2.8 93 2.8 105 ;
 END
END C PIN D DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 64.4 93 64.4 105 ;
 END
END D PIN E DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 198.8 39 198.8 39 ;
 END
END E PIN F DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 198.8 45 198.8 45 ;
 END
END F PIN G DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 2.8 111 2.8 111 ;
 END
END G
PIN VDD #here in the original was the pin declaratio missing!!!
PORT LAYER M2 ;
 WIDTH 3.6 ;
 PATH 1.8 27 199.8 27 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 PORT LAYER M2 ;
 WIDTH 3.6 ;
 PATH 1.8 57 199.8 57 ;
 END
END VSS OBS LAYER M2 ;
 RECT 1.0 80 66.2 166.5 ;
 RECT 1.0 1.5 200.6 23 ;
 RECT 1.0 31 200.6 53 ;
 RECT 1.0 61 200.6 82.5 ;
 # rectilinear shape description LAYER OVERLAP ;
 RECT 0 0 201.6 84 ;
 RECT 0 84 67.2 168 ;
 END
END LBLOCK

END LIBRARY
