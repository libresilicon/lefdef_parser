VIA VIABIGPOWER12 LAYER M1 ;
 RECT -21.0 -21.0 21.0 21.0 ;
 LAYER CUT12 ;
 RECT -2.4 -0.8 2.4 0.8 ;
 RECT -19.0 -19.0 -14.2 -17.4 ;
 RECT -19.0 17.4 -14.2 19.0;
 RECT 14.2 -19.0 19.0 -17.4 ;
 RECT 14.2 17.4 19.0 19.0 ;
 RECT -19.0 -0.8 -14.2 0.8 ;
 RECT -2.4 -19.0 2.4 -17.4 ;
 RECT 14.2 -0.8 19 0.8 ;
 RECT -2.4 17.4 2.4 19.0 ;
 LAYER M2 ;
 RECT -21.0 -21.0 21.0 21.0 ;
END VIABIGPOWER12 
