MACRO AND2J
 EEQ AND2 ;
 FOREIGN AND2SJ ;
 SIZE 67.2 BY 48 ;
 SYMMETRY X Y ;
 ORIGIN 0 6 ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 33 42 33 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 42 15 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 42 3 ;
 END
END B PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 -1.4 50.4 37.4 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 -1.4 16.8 37.4 ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 34.5 ;
 END
END AND2J 
