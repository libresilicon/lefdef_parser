VIA VIACENTER12 LAYER M1 ;
 RECT -4.6 -2.2 4.6 2.2 ;
 LAYER CUT12 ;
 RECT -3.1 -0.8 -1.9 0.8 ;
 RECT 1.9 -0.8 3.1 0.8 ;
 LAYER M2 ;
 RECT -4.4 -2.0 4.4 2.0 ;
END VIACENTER12 
