MACRO OR2
 FOREIGN OR2S ;
 SIZE 67.2 BY 42 ;
 SYMMETRY X Y ;
 SITE CORE1 ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 25.2 39 42 39 ;
 END
END Z PIN A DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 15 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 25.2 3 ;
 END
END B PIN VDD DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 50.4 4.6 50.4 10.0 ;
 PATH 50.4 27.4 50.4 37.4 ;
 VIA 50.4 3 C2PW ;
 VIA 50.4 21 C2PW ;
 VIA 50.4 33 C2PW ;
 VIA 50.4 39 C2PW ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE FEEDTHRU ;
 PORT LAYER M1 ;
 WIDTH 5.6 ;
 PATH 16.8 4.6 16.8 10.0 ;
 PATH 16.8 27.4 16.8 37.4 ;
 VIA 16.8 3 C2NW ;
 VIA 16.8 15 C2NW ;
 VIA 16.8 21 C2NW ;
 VIA 16.8 33 C2NW ;
 VIA 16.8 39 C2NW ;
 END
END VSS OBS LAYER M1 ;
 RECT 24.1 1.5 43.5 40.5 ;
 END
END OR2
