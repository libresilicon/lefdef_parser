LAYER metal1
  TYPE			ROUTING ;
  DIRECTION		HORIZONTAL ;
  PITCH			0.200 ;
  OFFSET		0.000 ;
  PROPERTY LEF57_MINSTEP "MINSTEP 0.100 MAXEDGES 1 ;" ;
  WIDTH			0.100 ;
  MAXWIDTH		10.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.40    0.46    1.40    4.10
  WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
  WIDTH    0.30         0.10    0.12    0.12    0.12    0.12
  WIDTH    0.46         0.10    0.12    0.15    0.15    0.15
  WIDTH    1.40         0.10    0.12    0.15    0.52    0.52
  WIDTH    4.10         0.10    0.12    0.15    0.52    1.40 ;

  PROPERTY LEF57_SPACING "SPACING 0.11 ENDOFLINE 0.12 WITHIN 0.045 PARALLELEDGE 0.11 WITHIN 0.11 ;" ;
  AREA 			0.041 ;
  MINENCLOSEDAREA	0.30 ;

  MINIMUMCUT 2 WIDTH 0.400 ;
  MINIMUMCUT 4 WIDTH 0.720 ;
  MINIMUMCUT 2 WIDTH 0.400 LENGTH 0.400 WITHIN 0.820 ;
  MINIMUMCUT 2 WIDTH 2.100 LENGTH 2.100 WITHIN 2.100 ;
  MINIMUMCUT 2 WIDTH 3.200 LENGTH 8.000 WITHIN 5.200 ;

END metal1
