MACRO IN1X
 class pad ;
 FOREIGN IN1X ;
 SIZE 151.2 BY 444 ;
 SYMMETRY X ;
 SITE IOX ;
 PIN Z DIRECTION OUTPUT ;
   PORT
   LAYER M1 ;
      PATH 61.6 444 72.8 444 ;
   END
 END Z
PIN PO
   DIRECTION OUTPUT ;
   PORT
     LAYER M1 ;
     PATH 78.4 444 84.0 444 ;
   END
  END PO
  PIN A
   DIRECTION INPUT ;
   PORT
      LAYER M1 ;
      PATH 95.2 444 100.8 444 ;
   END
   END A
  PIN PI
   DIRECTION INPUT ;
   PORT
   LAYER M1 ;
   PATH 106.4 444 112 444 ;
  END
 END PI
 PIN VDD
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      WIDTH 20 ;
      PATH 10 200 141.2 200 ;
    END
 END VDD
 PIN VSS
 DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT
   LAYER M1 ;
   WIDTH 20 ;
   PATH 10 100 141.2 100 ;
 END
END VSS
END IN1X 
