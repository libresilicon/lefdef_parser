MACRO LBLOCK
 FOREIGN LBLOCKS ;
 CLASS RING ;
 SIZE 201.6 BY 168 ;
 SITE LBLOCK ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 2.8 15 198.8 15 ;
 END
END Z PIN A DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 2.8 81 137.2 81 ;
 PATH 137.2 81 137.2 69 ;
 PATH 137.2 69 198.8 69 ;
 END
END A
PIN B DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 2.8 165 64.4 165 ;
 END
END B PIN C DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 2.8 93 2.8 105 ;
 END
END C PIN D DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 64.4 93 64.4 105 ;
 END
END D PIN E DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 198.8 39 198.8 39 ;
 END
END E PIN F DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 198.8 45 198.8 45 ;
 END
END F PIN G DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 2.8 111 2.8 111 ;
 END
END G
PIN VDD
 PORT LAYER M2 ;
 WIDTH 3.6 ;
 PATH 1.8 27 199.8 27 ;
 END
END VDD

PIN VSS DIRECTION INOUT ;
 PORT LAYER M2 ;
 WIDTH 3.6 ;
 PATH 1.8 57 199.8 57 ;
 END
END VSS OBS LAYER M2 ;
 RECT 1.0 80 66.2 166.5 ;
 RECT 1.0 1.5 200.6 23 ;
 RECT 1.0 31 200.6 53 ;
 RECT 1.0 61 200.6 82.5 ;
 # rectilinear shape description LAYER OVERLAP ;
 RECT 0 0 201.6 84 ;
 RECT 0 84 67.2 168 ;
 END
END LBLOCK
