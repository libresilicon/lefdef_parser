VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO h5
   CLASS BLOCK ;
   FOREIGN h5 ;
   ORIGIN 0 0 ;
   SIZE 303.2 BY 144 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1102_rst
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.19 0 284.29 0.51 ;
      END
   END FE_OFN1102_rst

   PIN FE_OFN267_n_4280
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.54 143.745 248.74 144 ;
      END
   END FE_OFN267_n_4280

   PIN FE_OFN827_n_3772
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 139.95 303.2 140.05 ;
      END
   END FE_OFN827_n_3772

   PIN FE_OFN829_n_8424
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.59 143.49 275.69 144 ;
      END
   END FE_OFN829_n_8424

   PIN n_10129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.75 0.51 120.85 ;
      END
   END n_10129

   PIN n_10572
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.95 0.51 136.05 ;
      END
   END n_10572

   PIN n_10650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.39 0 116.49 0.51 ;
      END
   END n_10650

   PIN n_10952
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.59 0 93.69 0.51 ;
      END
   END n_10952

   PIN n_10953
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.59 0 86.69 0.51 ;
      END
   END n_10953

   PIN n_12076
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.39 143.49 88.49 144 ;
      END
   END n_12076

   PIN n_12100
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.19 0 99.29 0.51 ;
      END
   END n_12100

   PIN n_12221
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.99 0 109.09 0.51 ;
      END
   END n_12221

   PIN n_1247
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 246.99 143.49 247.09 144 ;
      END
   END n_1247

   PIN n_12608
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.95 0.51 86.05 ;
      END
   END n_12608

   PIN n_12826
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.39 143.49 92.49 144 ;
      END
   END n_12826

   PIN n_13290
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.39 0 34.49 0.51 ;
      END
   END n_13290

   PIN n_13898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.35 0.51 85.45 ;
      END
   END n_13898

   PIN n_14243
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.39 0 86.49 0.51 ;
      END
   END n_14243

   PIN n_14244
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.59 0 92.69 0.51 ;
      END
   END n_14244

   PIN n_14522
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 253.99 143.49 254.09 144 ;
      END
   END n_14522

   PIN n_14855
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.59 0 104.69 0.51 ;
      END
   END n_14855

   PIN n_14856
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.39 0 104.49 0.51 ;
      END
   END n_14856

   PIN n_1487
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 71.55 303.2 71.65 ;
      END
   END n_1487

   PIN n_15005
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 120.15 303.2 120.25 ;
      END
   END n_15005

   PIN n_15031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.79 0 77.89 0.51 ;
      END
   END n_15031

   PIN n_15092
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.19 0 86.29 0.51 ;
      END
   END n_15092

   PIN n_15377
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 95.39 0 95.49 0.51 ;
      END
   END n_15377

   PIN n_1591
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.79 143.49 266.89 144 ;
      END
   END n_1591

   PIN n_15967
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 112.55 303.2 112.65 ;
      END
   END n_15967

   PIN n_16054
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.39 0 81.49 0.51 ;
      END
   END n_16054

   PIN n_16555
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.15 0.51 71.25 ;
      END
   END n_16555

   PIN n_16749
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.35 0.51 71.45 ;
      END
   END n_16749

   PIN n_16770
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.59 0 81.69 0.51 ;
      END
   END n_16770

   PIN n_17130
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.79 0 53.89 0.51 ;
      END
   END n_17130

   PIN n_17673
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.19 0 88.29 0.51 ;
      END
   END n_17673

   PIN n_19031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.15 0.51 76.25 ;
      END
   END n_19031

   PIN n_19333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.39 0 46.49 0.51 ;
      END
   END n_19333

   PIN n_19372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.75 0.51 71.85 ;
      END
   END n_19372

   PIN n_20390
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 13.55 303.2 13.65 ;
      END
   END n_20390

   PIN n_2339
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.79 143.49 48.89 144 ;
      END
   END n_2339

   PIN n_23513
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 40.35 303.2 40.45 ;
      END
   END n_23513

   PIN n_24465
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 225.79 0 225.89 0.51 ;
      END
   END n_24465

   PIN n_25465
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 228.39 143.49 228.49 144 ;
      END
   END n_25465

   PIN n_26031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 219.79 143.49 219.89 144 ;
      END
   END n_26031

   PIN n_27335
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 8.55 303.2 8.65 ;
      END
   END n_27335

   PIN n_28336
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 40.15 303.2 40.25 ;
      END
   END n_28336

   PIN n_28551
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.99 143.49 152.09 144 ;
      END
   END n_28551

   PIN n_28552
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.79 143.49 151.89 144 ;
      END
   END n_28552

   PIN n_28705
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 8.35 303.2 8.45 ;
      END
   END n_28705

   PIN n_29060
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 13.75 303.2 13.85 ;
      END
   END n_29060

   PIN n_29114
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.39 143.49 266.49 144 ;
      END
   END n_29114

   PIN n_29356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 119.95 303.2 120.05 ;
      END
   END n_29356

   PIN n_29588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 229.59 143.49 229.69 144 ;
      END
   END n_29588

   PIN n_29605
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 239.79 143.49 239.89 144 ;
      END
   END n_29605

   PIN n_2970
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.39 143.49 68.49 144 ;
      END
   END n_2970

   PIN n_3176
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 135.95 303.2 136.05 ;
      END
   END n_3176

   PIN n_3798
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.59 143.49 68.69 144 ;
      END
   END n_3798

   PIN n_3802
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.79 143.49 68.89 144 ;
      END
   END n_3802

   PIN n_3839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.39 143.49 50.49 144 ;
      END
   END n_3839

   PIN n_4058
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.39 143.49 59.49 144 ;
      END
   END n_4058

   PIN n_4072
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.79 143.49 80.89 144 ;
      END
   END n_4072

   PIN n_5262
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.59 143.49 266.69 144 ;
      END
   END n_5262

   PIN n_5327
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.19 143.49 266.29 144 ;
      END
   END n_5327

   PIN n_5340
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.99 143.49 52.09 144 ;
      END
   END n_5340

   PIN n_5341
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.59 143.49 41.69 144 ;
      END
   END n_5341

   PIN n_5519
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.39 143.49 248.49 144 ;
      END
   END n_5519

   PIN n_6244
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 94.75 0.51 94.85 ;
      END
   END n_6244

   PIN n_6256
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.99 143.49 78.09 144 ;
      END
   END n_6256

   PIN n_6595
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.59 0 103.69 0.51 ;
      END
   END n_6595

   PIN n_6979
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 94.35 0.51 94.45 ;
      END
   END n_6979

   PIN n_6987
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 94.55 0.51 94.65 ;
      END
   END n_6987

   PIN n_7017
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.59 143.49 5.69 144 ;
      END
   END n_7017

   PIN n_7224
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 122.59 143.49 122.69 144 ;
      END
   END n_7224

   PIN n_7237
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 94.55 303.2 94.65 ;
      END
   END n_7237

   PIN n_7274
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.39 143.49 61.49 144 ;
      END
   END n_7274

   PIN n_7311
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 239.59 143.49 239.69 144 ;
      END
   END n_7311

   PIN n_8443
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.19 143.49 80.29 144 ;
      END
   END n_8443

   PIN n_8444
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.59 143.49 77.69 144 ;
      END
   END n_8444

   PIN n_9230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.35 0.51 107.45 ;
      END
   END n_9230

   PIN n_9350
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.15 0.51 120.25 ;
      END
   END n_9350

   PIN n_9351
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.35 0.51 120.45 ;
      END
   END n_9351

   PIN n_9728
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.55 0.51 85.65 ;
      END
   END n_9728

   PIN n_9943
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.19 143.49 116.29 144 ;
      END
   END n_9943

   PIN x_out_21_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 76.35 303.2 76.45 ;
      END
   END x_out_21_1

   PIN x_out_21_22
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 112.35 303.2 112.45 ;
      END
   END x_out_21_22

   PIN x_out_21_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 67.35 303.2 67.45 ;
      END
   END x_out_21_23

   PIN x_out_21_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 121.55 303.2 121.65 ;
      END
   END x_out_21_24

   PIN x_out_21_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 93.95 303.2 94.05 ;
      END
   END x_out_21_25

   PIN x_out_21_26
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 62.15 303.2 62.25 ;
      END
   END x_out_21_26

   PIN x_out_25_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 40.55 303.2 40.65 ;
      END
   END x_out_25_29

   PIN x_out_25_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 22.35 303.2 22.45 ;
      END
   END x_out_25_30

   PIN x_out_53_22
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 84.95 303.2 85.05 ;
      END
   END x_out_53_22

   PIN x_out_53_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 112.35 303.2 112.45 ;
      END
   END x_out_53_24

   PIN x_out_53_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 94.35 303.2 94.45 ;
      END
   END x_out_53_25

   PIN x_out_53_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 112.15 303.2 112.25 ;
      END
   END x_out_53_28

   PIN x_out_55_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 121.35 303.2 121.45 ;
      END
   END x_out_55_14

   PIN x_out_57_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 93.55 303.2 93.65 ;
      END
   END x_out_57_29

   PIN x_out_57_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 84.75 303.2 84.85 ;
      END
   END x_out_57_30

   PIN x_out_5_13
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 104.15 303.2 104.25 ;
      END
   END x_out_5_13

   PIN FE_OFN1171_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.99 0 292.09 0.51 ;
      END
   END FE_OFN1171_n_4860

   PIN FE_OFN1264_n_29354
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.59 143.49 284.69 144 ;
      END
   END FE_OFN1264_n_29354

   PIN FE_OFN184_n_29402
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 103.95 303.2 104.05 ;
      END
   END FE_OFN184_n_29402

   PIN FE_OFN248_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.945 84.3 303.2 84.5 ;
      END
   END FE_OFN248_n_4162

   PIN FE_OFN261_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.39 143.49 96.49 144 ;
      END
   END FE_OFN261_n_4280

   PIN FE_OFN300_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 254.54 143.745 254.74 144 ;
      END
   END FE_OFN300_n_3069

   PIN FE_OFN303_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 243.14 0 243.34 0.255 ;
      END
   END FE_OFN303_n_3069

   PIN FE_OFN308_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.19 143.49 267.29 144 ;
      END
   END FE_OFN308_n_3069

   PIN FE_OFN326_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 239.54 143.745 239.74 144 ;
      END
   END FE_OFN326_n_4860

   PIN FE_OFN347_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.945 70.3 303.2 70.5 ;
      END
   END FE_OFN347_n_4860

   PIN FE_OFN35_n_15183
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 192.79 143.49 192.89 144 ;
      END
   END FE_OFN35_n_15183

   PIN FE_OFN400_n_28303
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 265.74 0 265.94 0.255 ;
      END
   END FE_OFN400_n_28303

   PIN FE_OFN56_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 104.1 0.255 104.3 ;
      END
   END FE_OFN56_n_27012

   PIN FE_OFN89_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 263.94 143.745 264.14 144 ;
      END
   END FE_OFN89_n_27449

   PIN FE_OFN90_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.945 104.9 303.2 105.1 ;
      END
   END FE_OFN90_n_27449

   PIN FE_OFN91_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 264.79 143.49 264.89 144 ;
      END
   END FE_OFN91_n_27449

   PIN FE_OFN92_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 284.74 143.745 284.94 144 ;
      END
   END FE_OFN92_n_27449

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.945 120.5 303.2 120.7 ;
      END
   END ispd_clk

   PIN n_10128
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.55 0.51 120.65 ;
      END
   END n_10128

   PIN n_14910
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.75 0.51 85.85 ;
      END
   END n_14910

   PIN n_15268
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 70.95 303.2 71.05 ;
      END
   END n_15268

   PIN n_15269
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 76.15 303.2 76.25 ;
      END
   END n_15269

   PIN n_15378
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.99 0 73.09 0.51 ;
      END
   END n_15378

   PIN n_15877
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.59 0 77.69 0.51 ;
      END
   END n_15877

   PIN n_15878
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.39 0 69.49 0.51 ;
      END
   END n_15878

   PIN n_15922
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 55.95 303.2 56.05 ;
      END
   END n_15922

   PIN n_17184
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 71.35 303.2 71.45 ;
      END
   END n_17184

   PIN n_17474
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.59 0 55.69 0.51 ;
      END
   END n_17474

   PIN n_17671
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.79 0 85.89 0.51 ;
      END
   END n_17671

   PIN n_17672
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.39 0 88.49 0.51 ;
      END
   END n_17672

   PIN n_19032
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.95 0.51 76.05 ;
      END
   END n_19032

   PIN n_21830
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.79 0 288.89 0.51 ;
      END
   END n_21830

   PIN n_22019
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 291.34 143.745 291.54 144 ;
      END
   END n_22019

   PIN n_22492
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 288.59 0 288.69 0.51 ;
      END
   END n_22492

   PIN n_23182
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.15 0.51 40.25 ;
      END
   END n_23182

   PIN n_2343
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 66.75 303.2 66.85 ;
      END
   END n_2343

   PIN n_237
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 56.15 303.2 56.25 ;
      END
   END n_237

   PIN n_23813
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 29.14 143.745 29.34 144 ;
      END
   END n_23813

   PIN n_24424
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.79 143.49 41.89 144 ;
      END
   END n_24424

   PIN n_24865
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.99 143.49 69.09 144 ;
      END
   END n_24865

   PIN n_26084
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.59 143.49 59.69 144 ;
      END
   END n_26084

   PIN n_26271
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.55 0.51 112.65 ;
      END
   END n_26271

   PIN n_26570
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.95 0.51 120.05 ;
      END
   END n_26570

   PIN n_27334
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 8.15 303.2 8.25 ;
      END
   END n_27334

   PIN n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 122.54 143.745 122.74 144 ;
      END
   END n_27449

   PIN n_28550
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 148.79 143.49 148.89 144 ;
      END
   END n_28550

   PIN n_28597
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.59 143.49 281.69 144 ;
      END
   END n_28597

   PIN n_29046
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128.14 143.745 128.34 144 ;
      END
   END n_29046

   PIN n_29068
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 99.39 143.49 99.49 144 ;
      END
   END n_29068

   PIN n_29126
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.19 143.49 79.29 144 ;
      END
   END n_29126

   PIN n_29261
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.945 104.5 303.2 104.7 ;
      END
   END n_29261

   PIN n_29664
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.34 143.745 41.54 144 ;
      END
   END n_29664

   PIN n_29683
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.945 139.5 303.2 139.7 ;
      END
   END n_29683

   PIN n_5003
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 239.19 143.49 239.29 144 ;
      END
   END n_5003

   PIN n_5445
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.19 143.49 79.29 144 ;
      END
   END n_5445

   PIN n_546
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.39 143.49 128.49 144 ;
      END
   END n_546

   PIN n_7214
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 61.95 303.2 62.05 ;
      END
   END n_7214

   PIN n_8671
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.19 143.49 52.29 144 ;
      END
   END n_8671

   PIN rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 284.34 143.745 284.54 144 ;
      END
   END rst

   PIN x_in_39_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 70.75 303.2 70.85 ;
      END
   END x_in_39_13

   PIN x_in_39_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 67.75 303.2 67.85 ;
      END
   END x_in_39_14

   PIN x_in_39_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 71.15 303.2 71.25 ;
      END
   END x_in_39_15

   PIN x_in_42_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.39 0 73.49 0.51 ;
      END
   END x_in_42_1

   PIN x_in_42_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 33.95 303.2 34.05 ;
      END
   END x_in_42_10

   PIN x_in_42_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 239.59 0 239.69 0.51 ;
      END
   END x_in_42_11

   PIN x_in_42_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 75.95 303.2 76.05 ;
      END
   END x_in_42_12

   PIN x_in_42_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 95.55 303.2 95.65 ;
      END
   END x_in_42_13

   PIN x_in_42_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 95.35 303.2 95.45 ;
      END
   END x_in_42_14

   PIN x_in_42_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 104.95 303.2 105.05 ;
      END
   END x_in_42_15

   PIN x_in_43_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 24.15 303.2 24.25 ;
      END
   END x_in_43_0

   PIN x_in_43_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 49.55 303.2 49.65 ;
      END
   END x_in_43_1

   PIN x_in_43_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 95.15 303.2 95.25 ;
      END
   END x_in_43_10

   PIN x_in_43_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 71.54 143.745 71.74 144 ;
      END
   END x_in_43_11

   PIN x_in_43_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 85.55 303.2 85.65 ;
      END
   END x_in_43_12

   PIN x_in_43_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 159.19 143.49 159.29 144 ;
      END
   END x_in_43_13

   PIN x_in_43_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 173.99 143.49 174.09 144 ;
      END
   END x_in_43_14

   PIN x_in_43_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 112.95 303.2 113.05 ;
      END
   END x_in_43_15

   PIN x_in_43_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 22.95 303.2 23.05 ;
      END
   END x_in_43_2

   PIN x_in_43_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 34.35 303.2 34.45 ;
      END
   END x_in_43_3

   PIN x_in_43_4
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 170.34 143.745 170.54 144 ;
      END
   END x_in_43_4

   PIN x_in_43_5
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.945 77.5 303.2 77.7 ;
      END
   END x_in_43_5

   PIN x_in_43_6
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 62.35 303.2 62.45 ;
      END
   END x_in_43_6

   PIN x_in_43_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.69 77.15 303.2 77.25 ;
      END
   END x_in_43_7

   PIN x_in_43_8
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 302.945 69.1 303.2 69.3 ;
      END
   END x_in_43_8

   PIN x_in_43_9
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.945 85.7 303.2 85.9 ;
      END
   END x_in_43_9

   PIN x_out_21_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.59 143.49 257.69 144 ;
      END
   END x_out_21_15

   PIN x_out_21_20
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.39 143.49 272.49 144 ;
      END
   END x_out_21_20

   PIN x_out_21_21
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 247.19 143.49 247.29 144 ;
      END
   END x_out_21_21

   PIN x_out_25_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 302.69 71.75 303.2 71.85 ;
      END
   END x_out_25_15

   PIN x_out_53_26
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.79 143.49 257.89 144 ;
      END
   END x_out_53_26

   PIN x_out_57_31
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.55 0.51 71.65 ;
      END
   END x_out_57_31

   OBS
      LAYER via4 ;
         RECT 0 0 303.2 144 ;
      LAYER via3 ;
         RECT 0 0 303.2 144 ;
      LAYER via2 ;
         RECT 0 0 303.2 144 ;
      LAYER via1 ;
         RECT 0 0 303.2 144 ;
      LAYER metal5 ;
         RECT 0 0 303.2 144 ;
      LAYER metal4 ;
         RECT 0 0 303.2 144 ;
      LAYER metal3 ;
         RECT 0 0 303.2 144 ;
      LAYER metal2 ;
         RECT 0 0 303.2 144 ;
      LAYER metal1 ;
         RECT 0 0 303.2 144 ;
   END
END h5

MACRO h4
   CLASS BLOCK ;
   FOREIGN h4 ;
   ORIGIN 0 0 ;
   SIZE 311 BY 212 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN276_n_16893
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.05 211.49 3.15 212 ;
      END
   END FE_OFN276_n_16893

   PIN FE_OFN282_n_7349
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 145.95 0.51 146.05 ;
      END
   END FE_OFN282_n_7349

   PIN FE_OFN339_n_4860
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 189.55 0.51 189.65 ;
      END
   END FE_OFN339_n_4860

   PIN FE_OFN352_n_4860
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 152.3 0.255 152.5 ;
      END
   END FE_OFN352_n_4860

   PIN n_10750
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.55 0.51 85.65 ;
      END
   END n_10750

   PIN n_12144
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.65 211.49 173.75 212 ;
      END
   END n_12144

   PIN n_1289
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.65 211.49 139.75 212 ;
      END
   END n_1289

   PIN n_13764
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 202.95 0.51 203.05 ;
      END
   END n_13764

   PIN n_14521
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.45 211.49 197.55 212 ;
      END
   END n_14521

   PIN n_14885
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 185.15 0.51 185.25 ;
      END
   END n_14885

   PIN n_15325
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.55 0.51 124.65 ;
      END
   END n_15325

   PIN n_15907
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.95 0.51 185.05 ;
      END
   END n_15907

   PIN n_16753
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.35 0.51 139.45 ;
      END
   END n_16753

   PIN n_16798
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 157.95 0.51 158.05 ;
      END
   END n_16798

   PIN n_17335
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 194.15 0.51 194.25 ;
      END
   END n_17335

   PIN n_17762
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.55 0.51 203.65 ;
      END
   END n_17762

   PIN n_17906
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.75 0.51 189.85 ;
      END
   END n_17906

   PIN n_17993
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 194.95 0.51 195.05 ;
      END
   END n_17993

   PIN n_18103
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.35 0.51 116.45 ;
      END
   END n_18103

   PIN n_18127
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.55 0.51 131.65 ;
      END
   END n_18127

   PIN n_18128
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.35 0.51 131.45 ;
      END
   END n_18128

   PIN n_18481
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.15 0.51 203.25 ;
      END
   END n_18481

   PIN n_18575
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.55 0.51 116.65 ;
      END
   END n_18575

   PIN n_1865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.25 211.49 123.35 212 ;
      END
   END n_1865

   PIN n_18833
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.75 0.51 131.85 ;
      END
   END n_18833

   PIN n_18835
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.15 0.51 131.25 ;
      END
   END n_18835

   PIN n_19121
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.55 0.51 189.65 ;
      END
   END n_19121

   PIN n_19140
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 202.95 0.51 203.05 ;
      END
   END n_19140

   PIN n_19235
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 194.75 0.51 194.85 ;
      END
   END n_19235

   PIN n_19322
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.15 0.51 87.25 ;
      END
   END n_19322

   PIN n_19382
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.35 0.51 58.45 ;
      END
   END n_19382

   PIN n_19891
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.55 0.51 139.65 ;
      END
   END n_19891

   PIN n_19966
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.35 0.51 203.45 ;
      END
   END n_19966

   PIN n_20233
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.95 0.51 140.05 ;
      END
   END n_20233

   PIN n_20283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 185.15 0.51 185.25 ;
      END
   END n_20283

   PIN n_20288
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.75 0.51 161.85 ;
      END
   END n_20288

   PIN n_20344
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.95 0.51 96.05 ;
      END
   END n_20344

   PIN n_20690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 203.15 0.51 203.25 ;
      END
   END n_20690

   PIN n_20766
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 175.35 0.51 175.45 ;
      END
   END n_20766

   PIN n_21207
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 202.75 0.51 202.85 ;
      END
   END n_21207

   PIN n_21332
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.75 0.51 85.85 ;
      END
   END n_21332

   PIN n_21382
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 45.45 211.49 45.55 212 ;
      END
   END n_21382

   PIN n_21383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.45 211.49 49.55 212 ;
      END
   END n_21383

   PIN n_21442
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 175.95 0.51 176.05 ;
      END
   END n_21442

   PIN n_21523
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.95 0.51 117.05 ;
      END
   END n_21523

   PIN n_22114
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.35 0.51 167.45 ;
      END
   END n_22114

   PIN n_22537
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.15 0.51 116.25 ;
      END
   END n_22537

   PIN n_22682
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.15 0.51 195.25 ;
      END
   END n_22682

   PIN n_22691
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.35 0.51 189.45 ;
      END
   END n_22691

   PIN n_22799
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.55 0.51 167.65 ;
      END
   END n_22799

   PIN n_23517
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.75 0.51 167.85 ;
      END
   END n_23517

   PIN n_23682
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.75 0.51 203.85 ;
      END
   END n_23682

   PIN n_23683
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 194.55 0.51 194.65 ;
      END
   END n_23683

   PIN n_23747
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.65 211.49 256.75 212 ;
      END
   END n_23747

   PIN n_23770
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.55 0.51 161.65 ;
      END
   END n_23770

   PIN n_23771
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.35 0.51 161.45 ;
      END
   END n_23771

   PIN n_24387
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.55 0.51 160.65 ;
      END
   END n_24387

   PIN n_24576
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.15 0.51 168.25 ;
      END
   END n_24576

   PIN n_25009
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 175.15 0.51 175.25 ;
      END
   END n_25009

   PIN n_25062
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 146.55 0.51 146.65 ;
      END
   END n_25062

   PIN n_25138
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 101.55 0.51 101.65 ;
      END
   END n_25138

   PIN n_2520
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 144.55 0.51 144.65 ;
      END
   END n_2520

   PIN n_2536
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 181.85 211.49 181.95 212 ;
      END
   END n_2536

   PIN n_25410
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.35 0.51 160.45 ;
      END
   END n_25410

   PIN n_25427
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 94.25 211.49 94.35 212 ;
      END
   END n_25427

   PIN n_26633
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 113.35 0.51 113.45 ;
      END
   END n_26633

   PIN n_27097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.05 211.49 114.15 212 ;
      END
   END n_27097

   PIN n_27589
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 114.05 211.49 114.15 212 ;
      END
   END n_27589

   PIN n_27724
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.75 0.51 116.85 ;
      END
   END n_27724

   PIN n_27869
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.65 211.49 290.75 212 ;
      END
   END n_27869

   PIN n_28230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 157.75 0.51 157.85 ;
      END
   END n_28230

   PIN n_28326
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.85 211.49 151.95 212 ;
      END
   END n_28326

   PIN n_28704
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 160.35 311 160.45 ;
      END
   END n_28704

   PIN n_28807
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.85 211.49 97.95 212 ;
      END
   END n_28807

   PIN n_28821
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 146.35 0.51 146.45 ;
      END
   END n_28821

   PIN n_29052
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.55 0.51 32.65 ;
      END
   END n_29052

   PIN n_29059
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 68.35 0.51 68.45 ;
      END
   END n_29059

   PIN n_29152
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.55 0.51 42.65 ;
      END
   END n_29152

   PIN n_29153
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.35 0.51 42.45 ;
      END
   END n_29153

   PIN n_29372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.75 0.51 32.85 ;
      END
   END n_29372

   PIN n_2947
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.35 0.51 72.45 ;
      END
   END n_2947

   PIN n_2951
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.95 0.51 141.05 ;
      END
   END n_2951

   PIN n_4021
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 144.75 0.51 144.85 ;
      END
   END n_4021

   PIN n_4881
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 188.75 0.51 188.85 ;
      END
   END n_4881

   PIN n_5362
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 72.15 0.51 72.25 ;
      END
   END n_5362

   PIN n_5669
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.75 0.51 139.85 ;
      END
   END n_5669

   PIN n_7328
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.05 211.49 141.15 212 ;
      END
   END n_7328

   PIN n_8581
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 113.55 0.51 113.65 ;
      END
   END n_8581

   PIN n_9651
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.95 0.51 68.05 ;
      END
   END n_9651

   PIN x_out_22_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 130.95 0.51 131.05 ;
      END
   END x_out_22_12

   PIN x_out_22_13
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 86.35 0.51 86.45 ;
      END
   END x_out_22_13

   PIN x_out_22_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 41.15 0.51 41.25 ;
      END
   END x_out_22_14

   PIN x_out_22_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.35 0.51 32.45 ;
      END
   END x_out_22_15

   PIN x_out_22_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 158.75 0.51 158.85 ;
      END
   END x_out_22_23

   PIN x_out_22_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 167.15 0.51 167.25 ;
      END
   END x_out_22_25

   PIN x_out_22_26
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 166.95 0.51 167.05 ;
      END
   END x_out_22_26

   PIN x_out_22_27
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 187.85 211.49 187.95 212 ;
      END
   END x_out_22_27

   PIN x_out_22_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.15 0.51 167.25 ;
      END
   END x_out_22_28

   PIN x_out_27_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 158.55 0.51 158.65 ;
      END
   END x_out_27_0

   PIN x_out_2_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 158.55 0.51 158.65 ;
      END
   END x_out_2_12

   PIN x_out_2_13
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.35 0.51 32.45 ;
      END
   END x_out_2_13

   PIN x_out_2_27
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 185.35 0.51 185.45 ;
      END
   END x_out_2_27

   PIN x_out_2_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 180.35 0.51 180.45 ;
      END
   END x_out_2_28

   PIN x_out_2_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 203.35 0.51 203.45 ;
      END
   END x_out_2_29

   PIN x_out_2_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 87.65 211.49 87.75 212 ;
      END
   END x_out_2_30

   PIN x_out_34_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 131.35 0.51 131.45 ;
      END
   END x_out_34_15

   PIN x_out_34_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 159.15 0.51 159.25 ;
      END
   END x_out_34_28

   PIN x_out_34_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 203.55 0.51 203.65 ;
      END
   END x_out_34_29

   PIN x_out_34_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.45 211.49 104.55 212 ;
      END
   END x_out_34_30

   PIN x_out_34_31
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 167.55 0.51 167.65 ;
      END
   END x_out_34_31

   PIN x_out_54_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 160.15 311 160.25 ;
      END
   END x_out_54_10

   PIN x_out_54_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 158.35 0.51 158.45 ;
      END
   END x_out_54_11

   PIN x_out_54_14
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 124.75 0.51 124.85 ;
      END
   END x_out_54_14

   PIN x_out_54_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.15 0.51 124.25 ;
      END
   END x_out_54_15

   PIN x_out_54_22
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 77.55 0.51 77.65 ;
      END
   END x_out_54_22

   PIN x_out_54_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 150.05 211.49 150.15 212 ;
      END
   END x_out_54_23

   PIN x_out_54_25
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 194.15 0.51 194.25 ;
      END
   END x_out_54_25

   PIN x_out_54_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 188.95 0.51 189.05 ;
      END
   END x_out_54_29

   PIN x_out_54_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 139.75 0.51 139.85 ;
      END
   END x_out_54_30

   PIN x_out_54_9
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 185.55 311 185.65 ;
      END
   END x_out_54_9

   PIN x_out_59_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 166.55 0.51 166.65 ;
      END
   END x_out_59_0

   PIN FE_OFN101_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 149.6 211.745 149.8 212 ;
      END
   END FE_OFN101_n_27449

   PIN FE_OFN105_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165 211.745 165.2 212 ;
      END
   END FE_OFN105_n_27449

   PIN FE_OFN1109_rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 125.6 211.745 125.8 212 ;
      END
   END FE_OFN1109_rst

   PIN FE_OFN1119_rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 148.8 211.745 149 212 ;
      END
   END FE_OFN1119_rst

   PIN FE_OFN133_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.5 0.255 188.7 ;
      END
   END FE_OFN133_n_27449

   PIN FE_OFN138_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 145.9 0.255 146.1 ;
      END
   END FE_OFN138_n_27449

   PIN FE_OFN175_n_26184
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.75 0.51 184.85 ;
      END
   END FE_OFN175_n_26184

   PIN FE_OFN183_n_29402
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 57.55 311 57.65 ;
      END
   END FE_OFN183_n_29402

   PIN FE_OFN212_n_29661
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.95 0.51 189.05 ;
      END
   END FE_OFN212_n_29661

   PIN FE_OFN214_n_29687
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 194.85 211.49 194.95 212 ;
      END
   END FE_OFN214_n_29687

   PIN FE_OFN234_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.8 211.745 125 212 ;
      END
   END FE_OFN234_n_4162

   PIN FE_OFN253_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.5 0.255 140.7 ;
      END
   END FE_OFN253_n_4280

   PIN FE_OFN257_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.745 130.9 311 131.1 ;
      END
   END FE_OFN257_n_4280

   PIN FE_OFN271_n_16028
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 253.25 211.49 253.35 212 ;
      END
   END FE_OFN271_n_16028

   PIN FE_OFN275_n_16893
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.75 0.51 130.85 ;
      END
   END FE_OFN275_n_16893

   PIN FE_OFN286_n_29266
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.05 211.49 105.15 212 ;
      END
   END FE_OFN286_n_29266

   PIN FE_OFN294_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.9 0.255 161.1 ;
      END
   END FE_OFN294_n_3069

   PIN FE_OFN331_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 174.95 0.51 175.05 ;
      END
   END FE_OFN331_n_4860

   PIN FE_OFN349_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 126 211.745 126.2 212 ;
      END
   END FE_OFN349_n_4860

   PIN FE_OFN37_n_17184
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 125.25 211.49 125.35 212 ;
      END
   END FE_OFN37_n_17184

   PIN FE_OFN404_n_28303
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 195.6 211.745 195.8 212 ;
      END
   END FE_OFN404_n_28303

   PIN FE_OFN68_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.745 87.3 311 87.5 ;
      END
   END FE_OFN68_n_27012

   PIN FE_OFN78_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 174.9 0.255 175.1 ;
      END
   END FE_OFN78_n_27012

   PIN FE_OFN7_n_28597
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.05 0 198.15 0.51 ;
      END
   END FE_OFN7_n_28597

   PIN FE_OFN95_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 136.8 0 137 0.255 ;
      END
   END FE_OFN95_n_27449

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.4 211.745 248.6 212 ;
      END
   END ispd_clk

   PIN n_1135
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 168.05 211.49 168.15 212 ;
      END
   END n_1135

   PIN n_11937
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.55 0.51 86.65 ;
      END
   END n_11937

   PIN n_12098
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.55 0.51 77.65 ;
      END
   END n_12098

   PIN n_12562
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.35 0.51 124.45 ;
      END
   END n_12562

   PIN n_13053
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.75 0.51 42.85 ;
      END
   END n_13053

   PIN n_13876
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 174.15 0.51 174.25 ;
      END
   END n_13876

   PIN n_14512
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.95 0.51 124.05 ;
      END
   END n_14512

   PIN n_14515
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 145.75 0.51 145.85 ;
      END
   END n_14515

   PIN n_14997
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 228.85 211.49 228.95 212 ;
      END
   END n_14997

   PIN n_15183
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.65 211.49 83.75 212 ;
      END
   END n_15183

   PIN n_16917
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.95 0.51 132.05 ;
      END
   END n_16917

   PIN n_17248
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.15 0.51 189.25 ;
      END
   END n_17248

   PIN n_1774
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.65 211.49 185.75 212 ;
      END
   END n_1774

   PIN n_18484
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 193.95 0.51 194.05 ;
      END
   END n_18484

   PIN n_18834
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.95 0.51 131.05 ;
      END
   END n_18834

   PIN n_20042
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.15 0.51 59.25 ;
      END
   END n_20042

   PIN n_20287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.55 0.51 184.65 ;
      END
   END n_20287

   PIN n_21013
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 117.15 0.51 117.25 ;
      END
   END n_21013

   PIN n_21076
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.1 0.255 86.3 ;
      END
   END n_21076

   PIN n_21471
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.55 0.51 72.65 ;
      END
   END n_21471

   PIN n_21988
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 202.3 0.255 202.5 ;
      END
   END n_21988

   PIN n_22184
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.15 0.51 96.25 ;
      END
   END n_22184

   PIN n_22202
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.15 0.51 102.25 ;
      END
   END n_22202

   PIN n_22681
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 194.75 0.51 194.85 ;
      END
   END n_22681

   PIN n_22758
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 87.15 0.51 87.25 ;
      END
   END n_22758

   PIN n_23465
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.95 0.51 87.05 ;
      END
   END n_23465

   PIN n_23509
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.85 211.49 248.95 212 ;
      END
   END n_23509

   PIN n_24114
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.75 0.51 86.85 ;
      END
   END n_24114

   PIN n_24126
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.75 0.51 57.85 ;
      END
   END n_24126

   PIN n_24135
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 101.75 0.51 101.85 ;
      END
   END n_24135

   PIN n_24421
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.25 211.49 279.35 212 ;
      END
   END n_24421

   PIN n_24716
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.95 0.51 59.05 ;
      END
   END n_24716

   PIN n_24799
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 263.45 211.49 263.55 212 ;
      END
   END n_24799

   PIN n_25130
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 263.05 211.49 263.15 212 ;
      END
   END n_25130

   PIN n_25150
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.15 0.51 58.25 ;
      END
   END n_25150

   PIN n_25188
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 167.55 311 167.65 ;
      END
   END n_25188

   PIN n_25502
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 265.65 211.49 265.75 212 ;
      END
   END n_25502

   PIN n_25659
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.15 0.51 27.25 ;
      END
   END n_25659

   PIN n_25660
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.35 0.51 27.45 ;
      END
   END n_25660

   PIN n_25661
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.75 0.51 27.85 ;
      END
   END n_25661

   PIN n_25854
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.95 0.51 54.05 ;
      END
   END n_25854

   PIN n_26081
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 252.05 211.49 252.15 212 ;
      END
   END n_26081

   PIN n_26139
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 160.55 311 160.65 ;
      END
   END n_26139

   PIN n_26416
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 151.95 311 152.05 ;
      END
   END n_26416

   PIN n_26568
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 195.05 211.49 195.15 212 ;
      END
   END n_26568

   PIN n_26827
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 159.35 0.51 159.45 ;
      END
   END n_26827

   PIN n_26857
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 116.15 311 116.25 ;
      END
   END n_26857

   PIN n_27121
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 158.15 311 158.25 ;
      END
   END n_27121

   PIN n_27307
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 131.55 0.51 131.65 ;
      END
   END n_27307

   PIN n_27331
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 189.35 0.51 189.45 ;
      END
   END n_27331

   PIN n_27332
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.05 211.49 305.15 212 ;
      END
   END n_27332

   PIN n_27415
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.85 211.49 216.95 212 ;
      END
   END n_27415

   PIN n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 174.8 211.745 175 212 ;
      END
   END n_27449

   PIN n_27488
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 240.05 211.49 240.15 212 ;
      END
   END n_27488

   PIN n_27709
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 231 0 231.2 0.255 ;
      END
   END n_27709

   PIN n_27914
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 158.95 0.51 159.05 ;
      END
   END n_27914

   PIN n_28602
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 130.65 211.49 130.75 212 ;
      END
   END n_28602

   PIN n_28607
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 245.6 211.745 245.8 212 ;
      END
   END n_28607

   PIN n_29033
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 69 0 69.2 0.255 ;
      END
   END n_29033

   PIN n_29046
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 174.2 211.745 174.4 212 ;
      END
   END n_29046

   PIN n_29104
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 105.6 211.745 105.8 212 ;
      END
   END n_29104

   PIN n_29683
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.7 0.255 87.9 ;
      END
   END n_29683

   PIN n_29687
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 298.05 211.49 298.15 212 ;
      END
   END n_29687

   PIN n_29691
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.8 0 125 0.255 ;
      END
   END n_29691

   PIN n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 240 211.745 240.2 212 ;
      END
   END n_4280

   PIN n_4687
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 130.75 0.51 130.85 ;
      END
   END n_4687

   PIN n_4811
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.15 0.51 72.25 ;
      END
   END n_4811

   PIN n_5360
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 57.35 0.51 57.45 ;
      END
   END n_5360

   PIN n_5402
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.75 0.51 72.85 ;
      END
   END n_5402

   PIN n_5677
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.85 211.49 159.95 212 ;
      END
   END n_5677

   PIN n_5983
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 54.15 0.51 54.25 ;
      END
   END n_5983

   PIN n_6742
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.05 211.49 123.15 212 ;
      END
   END n_6742

   PIN n_6849
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.15 0.51 140.25 ;
      END
   END n_6849

   PIN n_7229
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.05 211.49 177.15 212 ;
      END
   END n_7229

   PIN n_7287
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 158.85 211.49 158.95 212 ;
      END
   END n_7287

   PIN n_7289
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 158.65 211.49 158.75 212 ;
      END
   END n_7289

   PIN n_7402
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.85 211.49 176.95 212 ;
      END
   END n_7402

   PIN n_7417
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.65 211.49 159.75 212 ;
      END
   END n_7417

   PIN n_8331
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.55 0.51 57.65 ;
      END
   END n_8331

   PIN n_8423
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.05 211.49 150.15 212 ;
      END
   END n_8423

   PIN n_8513
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.65 211.49 176.75 212 ;
      END
   END n_8513

   PIN n_8772
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.05 211.49 178.15 212 ;
      END
   END n_8772

   PIN n_8915
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.35 0.51 77.45 ;
      END
   END n_8915

   PIN n_9113
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.35 0.51 57.45 ;
      END
   END n_9113

   PIN n_9336
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 101.95 0.51 102.05 ;
      END
   END n_9336

   PIN n_9650
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.95 0.51 58.05 ;
      END
   END n_9650

   PIN n_9936
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.75 0.51 58.85 ;
      END
   END n_9936

   PIN x_in_16_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.55 0.51 180.65 ;
      END
   END x_in_16_10

   PIN x_in_16_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 140.35 0.51 140.45 ;
      END
   END x_in_16_11

   PIN x_in_16_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 104.55 0.51 104.65 ;
      END
   END x_in_16_12

   PIN x_in_16_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 60.55 0.51 60.65 ;
      END
   END x_in_16_13

   PIN x_in_16_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 59.55 0.51 59.65 ;
      END
   END x_in_16_14

   PIN x_in_16_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.15 0.51 42.25 ;
      END
   END x_in_16_15

   PIN x_in_16_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.45 211.49 15.55 212 ;
      END
   END x_in_16_3

   PIN x_in_16_4
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.95 0.51 204.05 ;
      END
   END x_in_16_4

   PIN x_in_16_5
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.95 0.51 168.05 ;
      END
   END x_in_16_5

   PIN x_in_16_6
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.65 211.49 44.75 212 ;
      END
   END x_in_16_6

   PIN x_in_16_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 175.35 0.51 175.45 ;
      END
   END x_in_16_7

   PIN x_in_17_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.55 0.51 27.65 ;
      END
   END x_in_17_15

   PIN x_in_17_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.35 0.51 87.45 ;
      END
   END x_in_17_2

   PIN x_in_17_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 141.3 0.255 141.5 ;
      END
   END x_in_17_3

   PIN x_in_17_4
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 144.7 0.255 144.9 ;
      END
   END x_in_17_4

   PIN x_in_17_5
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 86.7 0.255 86.9 ;
      END
   END x_in_17_5

   PIN x_in_17_6
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 97.9 0.255 98.1 ;
      END
   END x_in_17_6

   PIN x_in_17_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.3 0.255 68.5 ;
      END
   END x_in_17_7

   PIN x_in_17_8
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 57.7 0.255 57.9 ;
      END
   END x_in_17_8

   PIN x_in_26_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.05 211.49 257.15 212 ;
      END
   END x_in_26_10

   PIN x_in_26_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 194.55 0.51 194.65 ;
      END
   END x_in_26_11

   PIN x_in_26_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 310.49 145.55 311 145.65 ;
      END
   END x_in_26_12

   PIN x_in_26_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 113.75 0.51 113.85 ;
      END
   END x_in_26_13

   PIN x_in_26_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.95 0.51 115.05 ;
      END
   END x_in_26_14

   PIN x_in_26_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 194.35 0.51 194.45 ;
      END
   END x_in_26_15

   PIN x_in_27_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.05 211.49 159.15 212 ;
      END
   END x_in_27_10

   PIN x_in_27_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 159 211.745 159.2 212 ;
      END
   END x_in_27_11

   PIN x_in_27_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.05 211.49 186.15 212 ;
      END
   END x_in_27_12

   PIN x_in_27_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.45 211.49 198.55 212 ;
      END
   END x_in_27_13

   PIN x_in_27_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.85 211.49 185.95 212 ;
      END
   END x_in_27_14

   PIN x_in_27_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 182.05 211.49 182.15 212 ;
      END
   END x_in_27_15

   PIN x_in_27_9
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 168.25 211.49 168.35 212 ;
      END
   END x_in_27_9

   PIN x_out_22_21
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.85 211.49 140.95 212 ;
      END
   END x_out_22_21

   PIN x_out_22_22
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 276.25 211.49 276.35 212 ;
      END
   END x_out_22_22

   PIN x_out_2_31
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 89.05 211.49 89.15 212 ;
      END
   END x_out_2_31

   PIN x_out_34_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.75 0.51 152.85 ;
      END
   END x_out_34_12

   OBS
      LAYER via4 ;
         RECT 0 0 311 212 ;
      LAYER via3 ;
         RECT 0 0 311 212 ;
      LAYER via2 ;
         RECT 0 0 311 212 ;
      LAYER via1 ;
         RECT 0 0 311 212 ;
      LAYER metal5 ;
         RECT 0 0 311 212 ;
      LAYER metal4 ;
         RECT 0 0 311 212 ;
      LAYER metal3 ;
         RECT 0 0 311 212 ;
      LAYER metal2 ;
         RECT 0 0 311 212 ;
      LAYER metal1 ;
         RECT 0 0 311 212 ;
   END
END h4

MACRO h3
   CLASS BLOCK ;
   FOREIGN h3 ;
   ORIGIN 0 0 ;
   SIZE 696.8 BY 172 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1143_n_27012
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 547 0 547.2 0.255 ;
      END
   END FE_OFN1143_n_27012

   PIN FE_OFN1193_n_12908
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 403.25 0 403.35 0.51 ;
      END
   END FE_OFN1193_n_12908

   PIN FE_OFN612_n_5698
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.45 171.49 160.55 172 ;
      END
   END FE_OFN612_n_5698

   PIN FE_OFN734_n_22952
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.35 0.51 96.45 ;
      END
   END FE_OFN734_n_22952

   PIN FE_OFN750_n_20252
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.45 0 133.55 0.51 ;
      END
   END FE_OFN750_n_20252

   PIN n_10335
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.25 0 43.35 0.51 ;
      END
   END n_10335

   PIN n_10432
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 389.65 0 389.75 0.51 ;
      END
   END n_10432

   PIN n_11256
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.85 171.49 107.95 172 ;
      END
   END n_11256

   PIN n_11262
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 42.55 696.8 42.65 ;
      END
   END n_11262

   PIN n_11285
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.45 171.49 124.55 172 ;
      END
   END n_11285

   PIN n_11526
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 691.25 0 691.35 0.51 ;
      END
   END n_11526

   PIN n_12365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 395.45 0 395.55 0.51 ;
      END
   END n_12365

   PIN n_12646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 86.15 696.8 86.25 ;
      END
   END n_12646

   PIN n_13045
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.05 171.49 124.15 172 ;
      END
   END n_13045

   PIN n_13066
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 25.25 0 25.35 0.51 ;
      END
   END n_13066

   PIN n_13175
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.85 0 16.95 0.51 ;
      END
   END n_13175

   PIN n_13229
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.05 171.49 160.15 172 ;
      END
   END n_13229

   PIN n_13260
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.05 171.49 178.15 172 ;
      END
   END n_13260

   PIN n_1333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.45 171.49 43.55 172 ;
      END
   END n_1333

   PIN n_13379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 664.25 0 664.35 0.51 ;
      END
   END n_13379

   PIN n_13564
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 481.45 0 481.55 0.51 ;
      END
   END n_13564

   PIN n_13965
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 385.05 0 385.15 0.51 ;
      END
   END n_13965

   PIN n_14028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 42.75 696.8 42.85 ;
      END
   END n_14028

   PIN n_14346
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 118.85 171.49 118.95 172 ;
      END
   END n_14346

   PIN n_14354
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 436.65 0 436.75 0.51 ;
      END
   END n_14354

   PIN n_14355
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 439.25 0 439.35 0.51 ;
      END
   END n_14355

   PIN n_14407
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.45 0 10.55 0.51 ;
      END
   END n_14407

   PIN n_14580
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 565.25 171.49 565.35 172 ;
      END
   END n_14580

   PIN n_14926
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 69.55 696.8 69.65 ;
      END
   END n_14926

   PIN n_14927
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 96.55 696.8 96.65 ;
      END
   END n_14927

   PIN n_15065
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 51.95 696.8 52.05 ;
      END
   END n_15065

   PIN n_15131
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.25 171.49 112.35 172 ;
      END
   END n_15131

   PIN n_15879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.45 0 16.55 0.51 ;
      END
   END n_15879

   PIN n_15880
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.45 0 7.55 0.51 ;
      END
   END n_15880

   PIN n_15991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 547.25 171.49 547.35 172 ;
      END
   END n_15991

   PIN n_16350
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 457.25 0 457.35 0.51 ;
      END
   END n_16350

   PIN n_16586
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 7.25 0 7.35 0.51 ;
      END
   END n_16586

   PIN n_16635
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 547.25 171.49 547.35 172 ;
      END
   END n_16635

   PIN n_16639
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 422.05 171.49 422.15 172 ;
      END
   END n_16639

   PIN n_16640
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 421.65 171.49 421.75 172 ;
      END
   END n_16640

   PIN n_16886
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 421.85 171.49 421.95 172 ;
      END
   END n_16886

   PIN n_17035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.55 0.51 69.65 ;
      END
   END n_17035

   PIN n_17253
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 141.55 696.8 141.65 ;
      END
   END n_17253

   PIN n_17495
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 412.25 171.49 412.35 172 ;
      END
   END n_17495

   PIN n_18101
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.75 0.51 12.85 ;
      END
   END n_18101

   PIN n_18104
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 123.55 696.8 123.65 ;
      END
   END n_18104

   PIN n_18396
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 394.05 0 394.15 0.51 ;
      END
   END n_18396

   PIN n_18435
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 141.75 696.8 141.85 ;
      END
   END n_18435

   PIN n_18488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 13.15 0.51 13.25 ;
      END
   END n_18488

   PIN n_18650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.65 0 26.75 0.51 ;
      END
   END n_18650

   PIN n_18683
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 395.25 0 395.35 0.51 ;
      END
   END n_18683

   PIN n_18728
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 655.25 171.49 655.35 172 ;
      END
   END n_18728

   PIN n_18812
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.95 0.51 52.05 ;
      END
   END n_18812

   PIN n_18882
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.15 0.51 86.25 ;
      END
   END n_18882

   PIN n_19039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.05 171.49 106.15 172 ;
      END
   END n_19039

   PIN n_19298
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 31.65 0 31.75 0.51 ;
      END
   END n_19298

   PIN n_19968
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.25 0 88.35 0.51 ;
      END
   END n_19968

   PIN n_20250
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.05 0 63.15 0.51 ;
      END
   END n_20250

   PIN n_20474
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 363.45 0 363.55 0.51 ;
      END
   END n_20474

   PIN n_20562
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 121.65 0 121.75 0.51 ;
      END
   END n_20562

   PIN n_20792
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.95 0.51 10.05 ;
      END
   END n_20792

   PIN n_20875
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 537.05 0 537.15 0.51 ;
      END
   END n_20875

   PIN n_21178
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.25 171.49 124.35 172 ;
      END
   END n_21178

   PIN n_21295
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.55 0.51 61.65 ;
      END
   END n_21295

   PIN n_21341
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 70.65 0 70.75 0.51 ;
      END
   END n_21341

   PIN n_21463
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.45 0 211.55 0.51 ;
      END
   END n_21463

   PIN n_21562
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 109.95 696.8 110.05 ;
      END
   END n_21562

   PIN n_21991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 520.45 171.49 520.55 172 ;
      END
   END n_21991

   PIN n_2220
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 628.25 0 628.35 0.51 ;
      END
   END n_2220

   PIN n_23291
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 138.6 0 138.8 0.255 ;
      END
   END n_23291

   PIN n_2342
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 601.25 0 601.35 0.51 ;
      END
   END n_2342

   PIN n_24279
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.35 0.51 12.45 ;
      END
   END n_24279

   PIN n_24915
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.05 0 258.15 0.51 ;
      END
   END n_24915

   PIN n_25379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.25 0 79.35 0.51 ;
      END
   END n_25379

   PIN n_25402
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.05 0 79.15 0.51 ;
      END
   END n_25402

   PIN n_25645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.45 0 165.55 0.51 ;
      END
   END n_25645

   PIN n_27432
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.45 0 115.55 0.51 ;
      END
   END n_27432

   PIN n_276
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.85 0 124.95 0.51 ;
      END
   END n_276

   PIN n_27650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 264.65 0 264.75 0.51 ;
      END
   END n_27650

   PIN n_27750
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.55 0.51 96.65 ;
      END
   END n_27750

   PIN n_28369
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.45 0 257.55 0.51 ;
      END
   END n_28369

   PIN n_3620
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.25 171.49 165.35 172 ;
      END
   END n_3620

   PIN n_3621
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 180.05 171.49 180.15 172 ;
      END
   END n_3621

   PIN n_3811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 601.45 0 601.55 0.51 ;
      END
   END n_3811

   PIN n_3847
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 590.45 0 590.55 0.51 ;
      END
   END n_3847

   PIN n_4099
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 384.05 0 384.15 0.51 ;
      END
   END n_4099

   PIN n_4578
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.45 0 43.55 0.51 ;
      END
   END n_4578

   PIN n_4928
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 374.05 0 374.15 0.51 ;
      END
   END n_4928

   PIN n_5156
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.65 0 36.75 0.51 ;
      END
   END n_5156

   PIN n_5158
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.05 0 34.15 0.51 ;
      END
   END n_5158

   PIN n_5537
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.85 171.49 119.95 172 ;
      END
   END n_5537

   PIN n_5556
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.65 171.49 160.75 172 ;
      END
   END n_5556

   PIN n_5557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.25 171.49 160.35 172 ;
      END
   END n_5557

   PIN n_5601
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 583.45 0 583.55 0.51 ;
      END
   END n_5601

   PIN n_5602
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 583.25 0 583.35 0.51 ;
      END
   END n_5602

   PIN n_5637
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 619.25 0 619.35 0.51 ;
      END
   END n_5637

   PIN n_5689
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 673.25 0 673.35 0.51 ;
      END
   END n_5689

   PIN n_5794
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 420.85 171.49 420.95 172 ;
      END
   END n_5794

   PIN n_5845
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.65 171.49 171.75 172 ;
      END
   END n_5845

   PIN n_5928
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 169.05 171.49 169.15 172 ;
      END
   END n_5928

   PIN n_6420
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 637.25 0 637.35 0.51 ;
      END
   END n_6420

   PIN n_6538
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.05 171.49 188.15 172 ;
      END
   END n_6538

   PIN n_6631
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 385.25 0 385.35 0.51 ;
      END
   END n_6631

   PIN n_6646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 421.05 171.49 421.15 172 ;
      END
   END n_6646

   PIN n_7384
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.25 0 25.35 0.51 ;
      END
   END n_7384

   PIN n_8420
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 566.45 0 566.55 0.51 ;
      END
   END n_8420

   PIN n_9616
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 646.45 0 646.55 0.51 ;
      END
   END n_9616

   PIN n_9619
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 341.05 0 341.15 0.51 ;
      END
   END n_9619

   PIN n_9640
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.65 171.49 124.75 172 ;
      END
   END n_9640

   PIN n_9641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.45 171.49 124.55 172 ;
      END
   END n_9641

   PIN n_9644
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.45 171.49 151.55 172 ;
      END
   END n_9644

   PIN n_9838
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 61.55 696.8 61.65 ;
      END
   END n_9838

   PIN n_9937
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 250.05 171.49 250.15 172 ;
      END
   END n_9937

   PIN n_999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.95 0.51 136.05 ;
      END
   END n_999

   PIN x_out_12_27
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 574.25 0 574.35 0.51 ;
      END
   END x_out_12_27

   PIN x_out_12_28
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 376.25 171.49 376.35 172 ;
      END
   END x_out_12_28

   PIN x_out_12_31
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 565.45 0 565.55 0.51 ;
      END
   END x_out_12_31

   PIN x_out_17_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.95 0.51 43.05 ;
      END
   END x_out_17_24

   PIN x_out_17_7
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 205.45 0 205.55 0.51 ;
      END
   END x_out_17_7

   PIN x_out_17_8
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 42.35 0.51 42.45 ;
      END
   END x_out_17_8

   PIN x_out_18_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 150.35 0.51 150.45 ;
      END
   END x_out_18_1

   PIN x_out_18_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 88.45 0 88.55 0.51 ;
      END
   END x_out_18_12

   PIN x_out_1_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.25 0 275.35 0.51 ;
      END
   END x_out_1_11

   PIN x_out_30_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 565.25 0 565.35 0.51 ;
      END
   END x_out_30_3

   PIN x_out_30_4
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 520.25 0 520.35 0.51 ;
      END
   END x_out_30_4

   PIN x_out_33_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 70.45 0 70.55 0.51 ;
      END
   END x_out_33_10

   PIN x_out_33_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 70.25 0 70.35 0.51 ;
      END
   END x_out_33_12

   PIN x_out_42_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 250.45 0 250.55 0.51 ;
      END
   END x_out_42_24

   PIN x_out_44_23
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 476.85 0 476.95 0.51 ;
      END
   END x_out_44_23

   PIN x_out_44_26
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 538.05 0 538.15 0.51 ;
      END
   END x_out_44_26

   PIN x_out_49_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 33.15 0.51 33.25 ;
      END
   END x_out_49_10

   PIN x_out_49_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 15.55 0.51 15.65 ;
      END
   END x_out_49_24

   PIN x_out_49_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 106.45 0 106.55 0.51 ;
      END
   END x_out_49_32

   PIN x_out_62_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 628.05 0 628.15 0.51 ;
      END
   END x_out_62_11

   PIN FE_OFN1123_rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 297 0 297.2 0.255 ;
      END
   END FE_OFN1123_rst

   PIN FE_OFN1124_rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 268 0 268.2 0.255 ;
      END
   END FE_OFN1124_rst

   PIN FE_OFN116_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 583.2 0 583.4 0.255 ;
      END
   END FE_OFN116_n_27449

   PIN FE_OFN1181_rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 602.2 171.745 602.4 172 ;
      END
   END FE_OFN1181_rst

   PIN FE_OFN129_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 529.2 0 529.4 0.255 ;
      END
   END FE_OFN129_n_27449

   PIN FE_OFN131_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 110.7 0.255 110.9 ;
      END
   END FE_OFN131_n_27449

   PIN FE_OFN139_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 119 0 119.2 0.255 ;
      END
   END FE_OFN139_n_27449

   PIN FE_OFN173_n_22948
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.25 0 133.35 0.51 ;
      END
   END FE_OFN173_n_22948

   PIN FE_OFN199_n_29637
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 547.45 0 547.55 0.51 ;
      END
   END FE_OFN199_n_29637

   PIN FE_OFN206_n_28771
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 531.85 171.49 531.95 172 ;
      END
   END FE_OFN206_n_28771

   PIN FE_OFN235_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 601.6 171.745 601.8 172 ;
      END
   END FE_OFN235_n_4162

   PIN FE_OFN23_n_26609
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.05 0 283.15 0.51 ;
      END
   END FE_OFN23_n_26609

   PIN FE_OFN244_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118.4 0 118.6 0.255 ;
      END
   END FE_OFN244_n_4162

   PIN FE_OFN254_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 205.8 0 206 0.255 ;
      END
   END FE_OFN254_n_4280

   PIN FE_OFN266_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 470 171.745 470.2 172 ;
      END
   END FE_OFN266_n_4280

   PIN FE_OFN280_n_16656
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 322.25 171.49 322.35 172 ;
      END
   END FE_OFN280_n_16656

   PIN FE_OFN296_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 257.2 171.745 257.4 172 ;
      END
   END FE_OFN296_n_3069

   PIN FE_OFN310_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 529 171.745 529.2 172 ;
      END
   END FE_OFN310_n_3069

   PIN FE_OFN313_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 106.8 0 107 0.255 ;
      END
   END FE_OFN313_n_3069

   PIN FE_OFN335_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 548 0 548.2 0.255 ;
      END
   END FE_OFN335_n_4860

   PIN FE_OFN361_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 252.2 171.745 252.4 172 ;
      END
   END FE_OFN361_n_4860

   PIN FE_OFN3_n_28682
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 99.65 0 99.75 0.51 ;
      END
   END FE_OFN3_n_28682

   PIN FE_OFN4_n_28682
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 569.65 0 569.75 0.51 ;
      END
   END FE_OFN4_n_28682

   PIN FE_OFN553_n_9468
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 466.25 0 466.35 0.51 ;
      END
   END FE_OFN553_n_9468

   PIN FE_OFN56_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 610.4 0 610.6 0.255 ;
      END
   END FE_OFN56_n_27012

   PIN FE_OFN63_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 517.6 0 517.8 0.255 ;
      END
   END FE_OFN63_n_27012

   PIN FE_OFN695_n_19853
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 150.55 696.8 150.65 ;
      END
   END FE_OFN695_n_19853

   PIN FE_OFN733_n_22952
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.45 0 97.55 0.51 ;
      END
   END FE_OFN733_n_22952

   PIN FE_OFN80_n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.2 0 124.4 0.255 ;
      END
   END FE_OFN80_n_27012

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 557 0 557.2 0.255 ;
      END
   END ispd_clk

   PIN n_10089
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 551.45 0 551.55 0.51 ;
      END
   END n_10089

   PIN n_10416
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 110.55 696.8 110.65 ;
      END
   END n_10416

   PIN n_10590
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.25 171.49 119.35 172 ;
      END
   END n_10590

   PIN n_10591
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.85 171.49 105.95 172 ;
      END
   END n_10591

   PIN n_10729
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 335.25 0 335.35 0.51 ;
      END
   END n_10729

   PIN n_10751
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.65 0 43.75 0.51 ;
      END
   END n_10751

   PIN n_11036
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.25 0 16.35 0.51 ;
      END
   END n_11036

   PIN n_11157
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.65 0 42.75 0.51 ;
      END
   END n_11157

   PIN n_11245
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.85 0 79.95 0.51 ;
      END
   END n_11245

   PIN n_11246
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.05 0 70.15 0.51 ;
      END
   END n_11246

   PIN n_11255
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.05 171.49 108.15 172 ;
      END
   END n_11255

   PIN n_11257
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.85 171.49 96.95 172 ;
      END
   END n_11257

   PIN n_11258
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.25 171.49 151.35 172 ;
      END
   END n_11258

   PIN n_11261
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 86.35 696.8 86.45 ;
      END
   END n_11261

   PIN n_11288
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.45 0 61.55 0.51 ;
      END
   END n_11288

   PIN n_11289
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.25 0 61.35 0.51 ;
      END
   END n_11289

   PIN n_11700
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 485.25 0 485.35 0.51 ;
      END
   END n_11700

   PIN n_11930
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 493.65 0 493.75 0.51 ;
      END
   END n_11930

   PIN n_12647
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 85.95 696.8 86.05 ;
      END
   END n_12647

   PIN n_12770
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.25 0 59.35 0.51 ;
      END
   END n_12770

   PIN n_12860
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.85 0 500.95 0.51 ;
      END
   END n_12860

   PIN n_12861
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.25 0 500.35 0.51 ;
      END
   END n_12861

   PIN n_13489
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 500.65 0 500.75 0.51 ;
      END
   END n_13489

   PIN n_13775
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 529.25 0 529.35 0.51 ;
      END
   END n_13775

   PIN n_15151
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.05 0 4.15 0.51 ;
      END
   END n_15151

   PIN n_15466
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 696.29 141.55 696.8 141.65 ;
      END
   END n_15466

   PIN n_15467
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 135.95 696.8 136.05 ;
      END
   END n_15467

   PIN n_15726
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 159.55 696.8 159.65 ;
      END
   END n_15726

   PIN n_15952
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.65 0 16.75 0.51 ;
      END
   END n_15952

   PIN n_16194
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 141.35 696.8 141.45 ;
      END
   END n_16194

   PIN n_16346
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 543.25 171.49 543.35 172 ;
      END
   END n_16346

   PIN n_16852
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.25 0 7.35 0.51 ;
      END
   END n_16852

   PIN n_17198
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 253.25 0 253.35 0.51 ;
      END
   END n_17198

   PIN n_17337
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.55 0.51 24.65 ;
      END
   END n_17337

   PIN n_17343
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 150.95 696.8 151.05 ;
      END
   END n_17343

   PIN n_17394
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.35 0.51 69.45 ;
      END
   END n_17394

   PIN n_17493
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 565.45 171.49 565.55 172 ;
      END
   END n_17493

   PIN n_17810
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 409.25 171.49 409.35 172 ;
      END
   END n_17810

   PIN n_17907
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.95 0.51 13.05 ;
      END
   END n_17907

   PIN n_18098
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 395.25 171.49 395.35 172 ;
      END
   END n_18098

   PIN n_18350
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.85 0 60.95 0.51 ;
      END
   END n_18350

   PIN n_18487
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.55 0.51 12.65 ;
      END
   END n_18487

   PIN n_18727
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 657.05 171.49 657.15 172 ;
      END
   END n_18727

   PIN n_1878
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 520.25 171.49 520.35 172 ;
      END
   END n_1878

   PIN n_18914
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.45 0 31.55 0.51 ;
      END
   END n_18914

   PIN n_18915
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.05 0 32.15 0.51 ;
      END
   END n_18915

   PIN n_19090
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 150.75 696.8 150.85 ;
      END
   END n_19090

   PIN n_19923
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.95 0.51 34.05 ;
      END
   END n_19923

   PIN n_20095
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.25 171.49 106.35 172 ;
      END
   END n_20095

   PIN n_20160
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 696.29 141.75 696.8 141.85 ;
      END
   END n_20160

   PIN n_20293
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 201.65 0 201.75 0.51 ;
      END
   END n_20293

   PIN n_20322
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.25 171.49 16.35 172 ;
      END
   END n_20322

   PIN n_20561
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 121.85 0 121.95 0.51 ;
      END
   END n_20561

   PIN n_20563
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 121.25 0 121.35 0.51 ;
      END
   END n_20563

   PIN n_20717
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.25 0 187.35 0.51 ;
      END
   END n_20717

   PIN n_20876
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 533.05 0 533.15 0.51 ;
      END
   END n_20876

   PIN n_20978
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.05 0 61.15 0.51 ;
      END
   END n_20978

   PIN n_21000
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.25 0 97.35 0.51 ;
      END
   END n_21000

   PIN n_22275
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.05 0 97.15 0.51 ;
      END
   END n_22275

   PIN n_24278
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 12.35 0.51 12.45 ;
      END
   END n_24278

   PIN n_24691
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.25 0 85.35 0.51 ;
      END
   END n_24691

   PIN n_24916
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.25 0 79.35 0.51 ;
      END
   END n_24916

   PIN n_25378
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.85 0 78.95 0.51 ;
      END
   END n_25378

   PIN n_25680
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 470.4 171.745 470.6 172 ;
      END
   END n_25680

   PIN n_25987
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.65 0 267.75 0.51 ;
      END
   END n_25987

   PIN n_26637
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.65 0 7.75 0.51 ;
      END
   END n_26637

   PIN n_2673
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 423.65 0 423.75 0.51 ;
      END
   END n_2673

   PIN n_2696
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 641.65 0 641.75 0.51 ;
      END
   END n_2696

   PIN n_27012
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 646.2 171.745 646.4 172 ;
      END
   END n_27012

   PIN n_27270
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.25 0 106.35 0.51 ;
      END
   END n_27270

   PIN n_27933
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 610 0 610.2 0.255 ;
      END
   END n_27933

   PIN n_28094
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.55 0.51 123.65 ;
      END
   END n_28094

   PIN n_28101
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 141.55 0.51 141.65 ;
      END
   END n_28101

   PIN n_28102
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.75 0.51 141.85 ;
      END
   END n_28102

   PIN n_28263
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.55 0.51 141.65 ;
      END
   END n_28263

   PIN n_28319
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.25 0 115.35 0.51 ;
      END
   END n_28319

   PIN n_28325
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.25 0 99.35 0.51 ;
      END
   END n_28325

   PIN n_28330
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 696.29 96.35 696.8 96.45 ;
      END
   END n_28330

   PIN n_2834
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 376.05 0 376.15 0.51 ;
      END
   END n_2834

   PIN n_28362
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.85 171.49 257.95 172 ;
      END
   END n_28362

   PIN n_29100
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.25 171.49 43.35 172 ;
      END
   END n_29100

   PIN n_3020
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.25 171.49 142.35 172 ;
      END
   END n_3020

   PIN n_3082
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.25 171.49 196.35 172 ;
      END
   END n_3082

   PIN n_3781
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.45 171.49 133.55 172 ;
      END
   END n_3781

   PIN n_3853
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 372.05 0 372.15 0.51 ;
      END
   END n_3853

   PIN n_4057
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 210.65 171.49 210.75 172 ;
      END
   END n_4057

   PIN n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 471.4 171.745 471.6 172 ;
      END
   END n_4162

   PIN n_4270
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 138.8 171.745 139 172 ;
      END
   END n_4270

   PIN n_4400
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.25 171.49 133.35 172 ;
      END
   END n_4400

   PIN n_4454
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.05 0 502.15 0.51 ;
      END
   END n_4454

   PIN n_4577
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.05 0 43.15 0.51 ;
      END
   END n_4577

   PIN n_4890
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 371.45 0 371.55 0.51 ;
      END
   END n_4890

   PIN n_4929
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 374.25 0 374.35 0.51 ;
      END
   END n_4929

   PIN n_5157
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.25 0 69.35 0.51 ;
      END
   END n_5157

   PIN n_5243
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.85 171.49 159.95 172 ;
      END
   END n_5243

   PIN n_5264
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 485.85 0 485.95 0.51 ;
      END
   END n_5264

   PIN n_5283
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 682.25 0 682.35 0.51 ;
      END
   END n_5283

   PIN n_5338
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.25 0 367.35 0.51 ;
      END
   END n_5338

   PIN n_5487
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.45 171.49 149.55 172 ;
      END
   END n_5487

   PIN n_5539
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.65 171.49 93.75 172 ;
      END
   END n_5539

   PIN n_5554
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 142.05 171.49 142.15 172 ;
      END
   END n_5554

   PIN n_5664
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 94.05 171.49 94.15 172 ;
      END
   END n_5664

   PIN n_5925
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 375.85 0 375.95 0.51 ;
      END
   END n_5925

   PIN n_5926
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.05 0 367.15 0.51 ;
      END
   END n_5926

   PIN n_6258
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.85 171.49 123.95 172 ;
      END
   END n_6258

   PIN n_6285
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 367.25 0 367.35 0.51 ;
      END
   END n_6285

   PIN n_6311
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 630.65 0 630.75 0.51 ;
      END
   END n_6311

   PIN n_7765
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 150.4 171.745 150.6 172 ;
      END
   END n_7765

   PIN n_7796
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.85 171.49 93.95 172 ;
      END
   END n_7796

   PIN n_7797
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.45 171.49 73.55 172 ;
      END
   END n_7797

   PIN n_7802
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.05 171.49 151.15 172 ;
      END
   END n_7802

   PIN n_7810
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 628.05 0 628.15 0.51 ;
      END
   END n_7810

   PIN n_7823
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.25 171.49 124.35 172 ;
      END
   END n_7823

   PIN n_8345
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 35.25 0 35.35 0.51 ;
      END
   END n_8345

   PIN n_8346
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.85 0 33.95 0.51 ;
      END
   END n_8346

   PIN n_8489
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.05 0 72.15 0.51 ;
      END
   END n_8489

   PIN n_8490
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.85 0 51.95 0.51 ;
      END
   END n_8490

   PIN n_8919
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 0 43.95 0.51 ;
      END
   END n_8919

   PIN n_8920
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.05 0 52.15 0.51 ;
      END
   END n_8920

   PIN n_9440
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 673.45 0 673.55 0.51 ;
      END
   END n_9440

   PIN n_9482
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 493.25 0 493.35 0.51 ;
      END
   END n_9482

   PIN n_9617
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 607.85 0 607.95 0.51 ;
      END
   END n_9617

   PIN n_9637
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.05 171.49 93.15 172 ;
      END
   END n_9637

   PIN n_9645
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.85 171.49 150.95 172 ;
      END
   END n_9645

   PIN n_9662
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.85 0 49.95 0.51 ;
      END
   END n_9662

   PIN n_9663
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.65 0 49.75 0.51 ;
      END
   END n_9663

   PIN n_9664
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.85 0 42.95 0.51 ;
      END
   END n_9664

   PIN n_9737
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 61.25 0 61.35 0.51 ;
      END
   END n_9737

   PIN n_9961
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.65 0 52.75 0.51 ;
      END
   END n_9961

   PIN x_in_13_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 406.65 0 406.75 0.51 ;
      END
   END x_in_13_10

   PIN x_in_13_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 423.4 0 423.6 0.255 ;
      END
   END x_in_13_11

   PIN x_in_13_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 385.25 0 385.35 0.51 ;
      END
   END x_in_13_12

   PIN x_in_13_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 412.45 0 412.55 0.51 ;
      END
   END x_in_13_13

   PIN x_in_13_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 403.45 0 403.55 0.51 ;
      END
   END x_in_13_14

   PIN x_in_13_9
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.45 0 502.55 0.51 ;
      END
   END x_in_13_9

   PIN x_in_19_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 97 171.745 97.2 172 ;
      END
   END x_in_19_10

   PIN x_in_19_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 151.2 171.745 151.4 172 ;
      END
   END x_in_19_11

   PIN x_in_19_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 169.8 171.745 170 172 ;
      END
   END x_in_19_12

   PIN x_in_19_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 169 171.745 169.2 172 ;
      END
   END x_in_19_13

   PIN x_in_19_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 180.45 171.49 180.55 172 ;
      END
   END x_in_19_14

   PIN x_in_19_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 169.45 171.49 169.55 172 ;
      END
   END x_in_19_15

   PIN x_in_19_9
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 137 171.745 137.2 172 ;
      END
   END x_in_19_9

   PIN x_in_30_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 520.45 0 520.55 0.51 ;
      END
   END x_in_30_2

   PIN x_in_34_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 42.55 0.51 42.65 ;
      END
   END x_in_34_7

   PIN x_in_35_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.2 0 52.4 0.255 ;
      END
   END x_in_35_1

   PIN x_in_51_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 619.4 0 619.6 0.255 ;
      END
   END x_in_51_11

   PIN x_in_51_12
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 645.8 0 646 0.255 ;
      END
   END x_in_51_12

   PIN x_in_51_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 628.45 0 628.55 0.51 ;
      END
   END x_in_51_13

   PIN x_in_51_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 619.05 0 619.15 0.51 ;
      END
   END x_in_51_14

   PIN x_in_51_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 646.25 0 646.35 0.51 ;
      END
   END x_in_51_15

   PIN x_out_12_26
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 457.45 0 457.55 0.51 ;
      END
   END x_out_12_26

   PIN x_out_49_30
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.65 0 258.75 0.51 ;
      END
   END x_out_49_30

   OBS
      LAYER via4 ;
         RECT 0 0 696.8 172 ;
      LAYER via3 ;
         RECT 0 0 696.8 172 ;
      LAYER via2 ;
         RECT 0 0 696.8 172 ;
      LAYER via1 ;
         RECT 0 0 696.8 172 ;
      LAYER metal5 ;
         RECT 0 0 696.8 172 ;
      LAYER metal4 ;
         RECT 0 0 696.8 172 ;
      LAYER metal3 ;
         RECT 0 0 696.8 172 ;
      LAYER metal2 ;
         RECT 0 0 696.8 172 ;
      LAYER metal1 ;
         RECT 0 0 696.8 172 ;
   END
END h3

MACRO h2
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 332.6 BY 254 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN953_n_13421
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.65 253.49 42.75 254 ;
      END
   END FE_OFN953_n_13421

   PIN n_10046
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 97.95 0.51 98.05 ;
      END
   END n_10046

   PIN n_10214
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END n_10214

   PIN n_1203
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.65 253.49 80.75 254 ;
      END
   END n_1203

   PIN n_12798
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.55 0.51 115.65 ;
      END
   END n_12798

   PIN n_13206
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.55 0.51 142.65 ;
      END
   END n_13206

   PIN n_13818
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.45 253.49 98.55 254 ;
      END
   END n_13818

   PIN n_14891
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 98.85 253.49 98.95 254 ;
      END
   END n_14891

   PIN n_15558
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 48.45 253.49 48.55 254 ;
      END
   END n_15558

   PIN n_19720
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 61.05 253.49 61.15 254 ;
      END
   END n_19720

   PIN n_21108
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.85 253.49 74.95 254 ;
      END
   END n_21108

   PIN n_21121
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.85 253.49 54.95 254 ;
      END
   END n_21121

   PIN n_23262
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.05 253.49 63.15 254 ;
      END
   END n_23262

   PIN n_23263
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.65 253.49 62.75 254 ;
      END
   END n_23263

   PIN n_23336
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.65 253.49 81.75 254 ;
      END
   END n_23336

   PIN n_24991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.85 253.49 62.95 254 ;
      END
   END n_24991

   PIN n_25847
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.65 253.49 107.75 254 ;
      END
   END n_25847

   PIN n_26581
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.25 253.49 98.35 254 ;
      END
   END n_26581

   PIN n_26926
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.05 253.49 100.15 254 ;
      END
   END n_26926

   PIN n_29040
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 187.55 0.51 187.65 ;
      END
   END n_29040

   PIN n_29135
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.25 253.49 104.35 254 ;
      END
   END n_29135

   PIN n_4730
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.95 0.51 161.05 ;
      END
   END n_4730

   PIN n_8503
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.75 0.51 160.85 ;
      END
   END n_8503

   PIN n_9692
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.65 253.49 40.75 254 ;
      END
   END n_9692

   PIN x_out_43_6
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.05 253.49 81.15 254 ;
      END
   END x_out_43_6

   PIN FE_OFN130_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.2 253.745 80.4 254 ;
      END
   END FE_OFN130_n_27449

   PIN FE_OFN259_n_4280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 62.6 253.745 62.8 254 ;
      END
   END FE_OFN259_n_4280

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.4 253.745 81.6 254 ;
      END
   END ispd_clk

   PIN n_10045
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.55 0.51 88.65 ;
      END
   END n_10045

   PIN n_10212
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.15 0.51 160.25 ;
      END
   END n_10212

   PIN n_10216
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 126.15 0.51 126.25 ;
      END
   END n_10216

   PIN n_10754
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.55 0.51 43.65 ;
      END
   END n_10754

   PIN n_11148
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 181.95 0.51 182.05 ;
      END
   END n_11148

   PIN n_12194
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.55 0.51 61.65 ;
      END
   END n_12194

   PIN n_12199
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.75 0.51 33.85 ;
      END
   END n_12199

   PIN n_12200
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.55 0.51 196.65 ;
      END
   END n_12200

   PIN n_12214
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.95 0.51 126.05 ;
      END
   END n_12214

   PIN n_13421
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.35 0.51 142.45 ;
      END
   END n_13421

   PIN n_19060
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.55 0.51 169.65 ;
      END
   END n_19060

   PIN n_20037
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.05 253.49 72.15 254 ;
      END
   END n_20037

   PIN n_22693
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.85 253.49 80.95 254 ;
      END
   END n_22693

   PIN n_23388
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.65 253.49 71.75 254 ;
      END
   END n_23388

   PIN n_24201
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 223.95 0.51 224.05 ;
      END
   END n_24201

   PIN n_24202
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.75 0.51 214.85 ;
      END
   END n_24202

   PIN n_24640
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.55 0.51 214.65 ;
      END
   END n_24640

   PIN n_25569
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.05 253.49 81.15 254 ;
      END
   END n_25569

   PIN n_26279
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.45 253.49 105.55 254 ;
      END
   END n_26279

   PIN n_27379
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.85 253.49 107.95 254 ;
      END
   END n_27379

   PIN n_27380
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.45 253.49 102.55 254 ;
      END
   END n_27380

   PIN n_28713
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.85 253.49 101.95 254 ;
      END
   END n_28713

   PIN n_28714
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.25 253.49 102.35 254 ;
      END
   END n_28714

   PIN n_4859
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.55 0.51 33.65 ;
      END
   END n_4859

   PIN n_6377
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.35 0.51 33.45 ;
      END
   END n_6377

   PIN n_6378
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.15 0.51 33.25 ;
      END
   END n_6378

   PIN n_8054
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.55 0.51 160.65 ;
      END
   END n_8054

   PIN n_8528
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.35 0.51 160.45 ;
      END
   END n_8528

   PIN n_8602
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.95 0.51 33.05 ;
      END
   END n_8602

   PIN x_in_52_13
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.05 253.49 108.15 254 ;
      END
   END x_in_52_13

   PIN x_in_52_6
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.05 253.49 72.15 254 ;
      END
   END x_in_52_6

   PIN x_out_43_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 89.45 253.49 89.55 254 ;
      END
   END x_out_43_7

   OBS
      LAYER via4 ;
         RECT 0 0 332.6 254 ;
      LAYER via3 ;
         RECT 0 0 332.6 254 ;
      LAYER via2 ;
         RECT 0 0 332.6 254 ;
      LAYER via1 ;
         RECT 0 0 332.6 254 ;
      LAYER metal5 ;
         RECT 0 0 332.6 254 ;
      LAYER metal4 ;
         RECT 0 0 332.6 254 ;
      LAYER metal3 ;
         RECT 0 0 332.6 254 ;
      LAYER metal2 ;
         RECT 0 0 332.6 254 ;
      LAYER metal1 ;
         RECT 0 0 332.6 254 ;
   END
END h2

MACRO h1
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 303.6 BY 172 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1036_n_26168
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.95 0.51 17.05 ;
      END
   END FE_OFN1036_n_26168

   PIN n_10017
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 170.85 0 170.95 0.51 ;
      END
   END n_10017

   PIN n_11653
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.05 171.49 39.15 172 ;
      END
   END n_11653

   PIN n_12968
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.85 0 116.95 0.51 ;
      END
   END n_12968

   PIN n_12983
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.85 0 14.95 0.51 ;
      END
   END n_12983

   PIN n_13860
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.05 0 171.15 0.51 ;
      END
   END n_13860

   PIN n_14132
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.45 0 179.55 0.51 ;
      END
   END n_14132

   PIN n_14219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.65 0 109.75 0.51 ;
      END
   END n_14219

   PIN n_14273
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.25 0 114.35 0.51 ;
      END
   END n_14273

   PIN n_1985
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.85 0 197.95 0.51 ;
      END
   END n_1985

   PIN n_21165
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.85 0 278.95 0.51 ;
      END
   END n_21165

   PIN n_23487
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 96.55 303.6 96.65 ;
      END
   END n_23487

   PIN n_24189
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 233.85 0 233.95 0.51 ;
      END
   END n_24189

   PIN n_24437
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 121.95 303.6 122.05 ;
      END
   END n_24437

   PIN n_2458
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 180.85 0 180.95 0.51 ;
      END
   END n_2458

   PIN n_3332
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.85 0 179.95 0.51 ;
      END
   END n_3332

   PIN n_4937
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.05 0 198.15 0.51 ;
      END
   END n_4937

   PIN n_5596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.05 0 155.15 0.51 ;
      END
   END n_5596

   PIN n_5761
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 251.85 0 251.95 0.51 ;
      END
   END n_5761

   PIN n_5771
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 242.85 0 242.95 0.51 ;
      END
   END n_5771

   PIN n_5839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.65 0 179.75 0.51 ;
      END
   END n_5839

   PIN n_6223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 158.05 0 158.15 0.51 ;
      END
   END n_6223

   PIN n_6579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.05 0 125.15 0.51 ;
      END
   END n_6579

   PIN n_6722
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 215.85 0 215.95 0.51 ;
      END
   END n_6722

   PIN n_7868
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.45 0 233.55 0.51 ;
      END
   END n_7868

   PIN n_7889
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.85 0 152.95 0.51 ;
      END
   END n_7889

   PIN n_8086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54.05 0 54.15 0.51 ;
      END
   END n_8086

   PIN n_8089
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.05 0 196.15 0.51 ;
      END
   END n_8089

   PIN n_8142
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 143.85 0 143.95 0.51 ;
      END
   END n_8142

   PIN n_8523
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.85 0 224.95 0.51 ;
      END
   END n_8523

   PIN n_8596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.05 0 135.15 0.51 ;
      END
   END n_8596

   PIN n_8597
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.85 0 134.95 0.51 ;
      END
   END n_8597

   PIN n_8601
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.85 0 161.95 0.51 ;
      END
   END n_8601

   PIN n_8972
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.85 0 98.95 0.51 ;
      END
   END n_8972

   PIN x_out_29_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 69.95 303.6 70.05 ;
      END
   END x_out_29_0

   PIN x_out_29_1
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.95 0.51 53.05 ;
      END
   END x_out_29_1

   PIN x_out_37_21
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 303.09 87.75 303.6 87.85 ;
      END
   END x_out_37_21

   PIN x_out_38_12
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 303.09 96.55 303.6 96.65 ;
      END
   END x_out_38_12

   PIN x_out_6_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 114.55 303.6 114.65 ;
      END
   END x_out_6_10

   PIN x_out_6_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 60.55 303.6 60.65 ;
      END
   END x_out_6_11

   PIN FE_OFN251_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 69 171.745 69.2 172 ;
      END
   END FE_OFN251_n_4162

   PIN FE_OFN306_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.9 0.255 123.1 ;
      END
   END FE_OFN306_n_3069

   PIN FE_OFN324_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.345 122.9 303.6 123.1 ;
      END
   END FE_OFN324_n_4860

   PIN FE_OFN330_n_4860
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 233.8 171.745 234 172 ;
      END
   END FE_OFN330_n_4860

   PIN FE_OFN393_n_14663
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.05 171.49 53.15 172 ;
      END
   END FE_OFN393_n_14663

   PIN FE_OFN662_n_27899
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 155.35 0.51 155.45 ;
      END
   END FE_OFN662_n_27899

   PIN FE_OFN810_n_12878
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 51.95 303.6 52.05 ;
      END
   END FE_OFN810_n_12878

   PIN FE_OFN93_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.1 0.255 52.3 ;
      END
   END FE_OFN93_n_27449

   PIN FE_OFN96_n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 154.3 0.255 154.5 ;
      END
   END FE_OFN96_n_27449

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.3 0.255 85.5 ;
      END
   END ispd_clk

   PIN n_10004
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 226.65 0 226.75 0.51 ;
      END
   END n_10004

   PIN n_12575
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.85 0 186.95 0.51 ;
      END
   END n_12575

   PIN n_13218
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.85 0 233.95 0.51 ;
      END
   END n_13218

   PIN n_13671
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.45 0 231.55 0.51 ;
      END
   END n_13671

   PIN n_13859
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 170.85 0 170.95 0.51 ;
      END
   END n_13859

   PIN n_14448
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.65 0 233.75 0.51 ;
      END
   END n_14448

   PIN n_14791
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.85 0 220.95 0.51 ;
      END
   END n_14791

   PIN n_17925
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.65 171.49 14.75 172 ;
      END
   END n_17925

   PIN n_21076
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.345 42.5 303.6 42.7 ;
      END
   END n_21076

   PIN n_21393
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.35 0.51 122.45 ;
      END
   END n_21393

   PIN n_21394
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.15 0.51 122.25 ;
      END
   END n_21394

   PIN n_21551
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 264.05 0 264.15 0.51 ;
      END
   END n_21551

   PIN n_23020
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.85 171.49 30.95 172 ;
      END
   END n_23020

   PIN n_2355
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.85 0 188.95 0.51 ;
      END
   END n_2355

   PIN n_24577
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 121.95 0.51 122.05 ;
      END
   END n_24577

   PIN n_25555
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.55 0.51 114.65 ;
      END
   END n_25555

   PIN n_25843
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 84.95 0.51 85.05 ;
      END
   END n_25843

   PIN n_26168
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 303.09 9.95 303.6 10.05 ;
      END
   END n_26168

   PIN n_26689
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.95 0.51 108.05 ;
      END
   END n_26689

   PIN n_28608
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 154.7 0.255 154.9 ;
      END
   END n_28608

   PIN n_2901
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 207.65 0 207.75 0.51 ;
      END
   END n_2901

   PIN n_4914
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 170.65 0 170.75 0.51 ;
      END
   END n_4914

   PIN n_5242
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 227.85 0 227.95 0.51 ;
      END
   END n_5242

   PIN n_5597
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 252.05 0 252.15 0.51 ;
      END
   END n_5597

   PIN n_5828
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.85 0 175.95 0.51 ;
      END
   END n_5828

   PIN n_7867
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 242.85 0 242.95 0.51 ;
      END
   END n_7867

   PIN n_8074
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 219.85 0 219.95 0.51 ;
      END
   END n_8074

   PIN n_8076
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.65 0 224.75 0.51 ;
      END
   END n_8076

   PIN n_8650
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.65 0 197.75 0.51 ;
      END
   END n_8650

   PIN n_8971
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.05 0 98.15 0.51 ;
      END
   END n_8971

   PIN n_9998
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.05 0 234.15 0.51 ;
      END
   END n_9998

   PIN n_9999
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 243.05 0 243.15 0.51 ;
      END
   END n_9999

   PIN x_in_46_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 303.09 69.75 303.6 69.85 ;
      END
   END x_in_46_0

   PIN x_in_61_5
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.8 0 153 0.255 ;
      END
   END x_in_61_5

   PIN x_in_61_6
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 135.4 0 135.6 0.255 ;
      END
   END x_in_61_6

   PIN x_in_61_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.6 0 186.8 0.255 ;
      END
   END x_in_61_7

   PIN x_in_61_8
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 208.2 0 208.4 0.255 ;
      END
   END x_in_61_8

   PIN x_in_61_9
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 215.8 0 216 0.255 ;
      END
   END x_in_61_9

   OBS
      LAYER via4 ;
         RECT 0 0 303.6 172 ;
      LAYER via3 ;
         RECT 0 0 303.6 172 ;
      LAYER via2 ;
         RECT 0 0 303.6 172 ;
      LAYER via1 ;
         RECT 0 0 303.6 172 ;
      LAYER metal5 ;
         RECT 0 0 303.6 172 ;
      LAYER metal4 ;
         RECT 0 0 303.6 172 ;
      LAYER metal3 ;
         RECT 0 0 303.6 172 ;
      LAYER metal2 ;
         RECT 0 0 303.6 172 ;
      LAYER metal1 ;
         RECT 0 0 303.6 172 ;
   END
END h1

MACRO h0
   CLASS BLOCK ;
   FOREIGN h0 ;
   ORIGIN 0 0 ;
   SIZE 329.6 BY 158 ;
   SYMMETRY X Y R90 ;
   PIN n_13301
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.85 0 171.95 0.51 ;
      END
   END n_13301

   PIN n_13302
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.85 0 159.95 0.51 ;
      END
   END n_13302

   PIN n_13303
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.05 0 160.15 0.51 ;
      END
   END n_13303

   PIN n_13488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.05 0 223.15 0.51 ;
      END
   END n_13488

   PIN n_14077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 247.85 0 247.95 0.51 ;
      END
   END n_14077

   PIN n_14078
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 241.05 0 241.15 0.51 ;
      END
   END n_14078

   PIN n_14581
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 241.05 0 241.15 0.51 ;
      END
   END n_14581

   PIN n_15640
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.05 0 124.15 0.51 ;
      END
   END n_15640

   PIN n_15661
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 214.05 0 214.15 0.51 ;
      END
   END n_15661

   PIN n_16544
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 242.65 0 242.75 0.51 ;
      END
   END n_16544

   PIN n_19438
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.09 22.745 329.6 22.845 ;
      END
   END n_19438

   PIN n_20533
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.09 80.145 329.6 80.245 ;
      END
   END n_20533

   PIN n_3465
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.25 0 56.35 0.51 ;
      END
   END n_3465

   PIN n_6033
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 95.05 0 95.15 0.51 ;
      END
   END n_6033

   PIN n_7083
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.05 0 79.15 0.51 ;
      END
   END n_7083

   PIN n_7084
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.25 0 79.35 0.51 ;
      END
   END n_7084

   PIN x_out_15_20
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 191.45 157.49 191.55 158 ;
      END
   END x_out_15_20

   PIN x_out_15_24
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.09 128.345 329.6 128.445 ;
      END
   END x_out_15_24

   PIN FE_OFN1111_rst
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.345 28.095 329.6 28.295 ;
      END
   END FE_OFN1111_rst

   PIN FE_OFN17_n_29617
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 27.745 0.51 27.845 ;
      END
   END FE_OFN17_n_29617

   PIN FE_OFN251_n_4162
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 313.2 0 313.4 0.255 ;
      END
   END FE_OFN251_n_4162

   PIN FE_OFN288_n_29266
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.65 0 270.75 0.51 ;
      END
   END FE_OFN288_n_29266

   PIN FE_OFN314_n_3069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 240.6 0 240.8 0.255 ;
      END
   END FE_OFN314_n_3069

   PIN FE_OFN409_n_28303
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 137.295 0.255 137.495 ;
      END
   END FE_OFN409_n_28303

   PIN FE_OFN660_n_19445
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 277.05 0 277.15 0.51 ;
      END
   END FE_OFN660_n_19445

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 134 0 134.2 0.255 ;
      END
   END ispd_clk

   PIN n_10314
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.85 0 96.95 0.51 ;
      END
   END n_10314

   PIN n_10315
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.05 0 115.15 0.51 ;
      END
   END n_10315

   PIN n_11856
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.85 0 266.95 0.51 ;
      END
   END n_11856

   PIN n_15273
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.05 0 196.15 0.51 ;
      END
   END n_15273

   PIN n_17533
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 312.85 0 312.95 0.51 ;
      END
   END n_17533

   PIN n_18413
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 240.85 0 240.95 0.51 ;
      END
   END n_18413

   PIN n_20363
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 312.85 0 312.95 0.51 ;
      END
   END n_20363

   PIN n_21988
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 324.2 0 324.4 0.255 ;
      END
   END n_21988

   PIN n_27449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.345 79.695 329.6 79.895 ;
      END
   END n_27449

   PIN n_3028
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.05 0 56.15 0.51 ;
      END
   END n_3028

   PIN n_3132
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.25 0 57.35 0.51 ;
      END
   END n_3132

   PIN n_3771
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.85 0 87.95 0.51 ;
      END
   END n_3771

   PIN n_4593
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.45 0 69.55 0.51 ;
      END
   END n_4593

   PIN n_4594
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.85 0 68.95 0.51 ;
      END
   END n_4594

   PIN n_4873
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.85 0 60.95 0.51 ;
      END
   END n_4873

   PIN n_5057
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.65 0 69.75 0.51 ;
      END
   END n_5057

   PIN n_5315
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.85 0 56.95 0.51 ;
      END
   END n_5315

   PIN n_6966
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.85 0 78.95 0.51 ;
      END
   END n_6966

   PIN n_7082
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.65 0 85.75 0.51 ;
      END
   END n_7082

   PIN n_871
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.09 27.745 329.6 27.845 ;
      END
   END n_871

   PIN x_in_25_4
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.8 0 79 0.255 ;
      END
   END x_in_25_4

   PIN x_in_25_5
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.8 0 57 0.255 ;
      END
   END x_in_25_5

   PIN x_in_25_6
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.2 0 96.4 0.255 ;
      END
   END x_in_25_6

   PIN x_in_25_7
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 9.6 0 9.8 0.255 ;
      END
   END x_in_25_7

   PIN x_out_38_4
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 329.09 65.345 329.6 65.445 ;
      END
   END x_out_38_4

   OBS
      LAYER via4 ;
         RECT 0 0 329.6 158 ;
      LAYER via3 ;
         RECT 0 0 329.6 158 ;
      LAYER via2 ;
         RECT 0 0 329.6 158 ;
      LAYER via1 ;
         RECT 0 0 329.6 158 ;
      LAYER metal5 ;
         RECT 0 0 329.6 158 ;
      LAYER metal4 ;
         RECT 0 0 329.6 158 ;
      LAYER metal3 ;
         RECT 0 0 329.6 158 ;
      LAYER metal2 ;
         RECT 0 0 329.6 158 ;
      LAYER metal1 ;
         RECT 0 0 329.6 158 ;
   END
END h0

MACRO ms00f80
   CLASS CORE ;
   FOREIGN ms00f80 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN ck
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END ck

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END d

END ms00f80

MACRO no02f01
   CLASS CORE ;
   FOREIGN no02f01 ;
   ORIGIN 0 0 ;
   SIZE 0.8 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

END no02f01

MACRO oa12f01
   CLASS CORE ;
   FOREIGN oa12f01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END oa12f01

MACRO in01f01
   CLASS CORE ;
   FOREIGN in01f01 ;
   ORIGIN 0 0 ;
   SIZE 0.4 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

END in01f01

MACRO na02f01
   CLASS CORE ;
   FOREIGN na02f01 ;
   ORIGIN 0 0 ;
   SIZE 0.8 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

END na02f01

MACRO oa22f01
   CLASS CORE ;
   FOREIGN oa22f01 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

END oa22f01

MACRO ao22s01
   CLASS CORE ;
   FOREIGN ao22s01 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

END ao22s01

MACRO ao12f01
   CLASS CORE ;
   FOREIGN ao12f01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END ao12f01

MACRO no03m01
   CLASS CORE ;
   FOREIGN no03m01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END no03m01

MACRO na03f01
   CLASS CORE ;
   FOREIGN na03f01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END na03f01

END LIBRARY
