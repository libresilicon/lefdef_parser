VIARULE VIAGEN23 GENERATE
 LAYER M2 ;
 ENCLOSURE 0.01 0.05 ;
 LAYER M3 ;
 ENCLOSURE 0.01 0.05 ;
 LAYER CUT23 ;
 RECT -0.06 -0.06 0.06 0.06 ;
 SPACING 0.14 BY 0.14 ;
END VIAGEN23 
