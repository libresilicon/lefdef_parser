MACRO IN1Y EEQ IN1X ;
 FOREIGN IN1Y ;
 class pad ;
 SIZE 436.8 BY 150 ;
 SYMMETRY Y ;
 SITE IOY ;
 PIN Z DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      PATH 0 69 0 75 ;
    END
 END Z
 PIN PO
    DIRECTION OUTPUT ;
    PORT
      LAYER M2 ;
      PATH 0 81 0 87 ;
    END
 END PO
 PIN A DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 51 0 57 ;
 END
END A PIN PI DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 0 39 0 45 ;
 END
END PI PIN VDD DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 236.8 10 236.8 140 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE ABUTMENT ;
 PORT LAYER M2 ;
 WIDTH 20 ;
 PATH 336.8 10 336.8 140 ;
 END
END VSS
END IN1Y 
