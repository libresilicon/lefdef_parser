VIA VIA23 DEFAULT LAYER M3 ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT23 ;
 RECT -0.8 -0.8 0.8 0.8 ;
 LAYER M2 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END VIA23 
