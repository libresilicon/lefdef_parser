LAYER via2
  TYPE CUT ;
  SPACING		0.10 ;
  SPACING		0.13 ADJACENTCUTS 3 WITHIN 0.15 ;
  PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
END via2
