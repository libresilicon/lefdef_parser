MACRO I2BLOCK FOREIGN I2BLOCKS ;
 CLASS RING ;
 SIZE 672 BY 504 ;
 SITE I2BLOCK ;
 PIN Z DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 22.8 21 649.2 21 ;
 END
END Z PIN A DIRECTION OUTPUT ;
 PORT LAYER M2 ;
 PATH 22.8 63 154.0 63 ;
 PATH 154.0 63 154.0 129;
 PATH 154.0 129 447.6 129 ;
 END
END A PIN B DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 137.2 423 447.6 423 ;
 END
END B PIN C DIRECTION INPUT ;
 PORT LAYER M2 ;
 PATH 204.4 165 271.6 165 ;
 END
END C PIN D DIRECTION INPUT ;
PORT LAYER M2 ;
 PATH 204.4 171 271.6 171 ;
 END
END D PIN E DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 204.4 213 204.4 213 ;
 END
END E PIN F DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 406 249 406 273 ;
 END
END F PIN G DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 338.8 249 338.8 273 ;
 END
END G PIN H DIRECTION INPUT ;
 PORT LAYER M1 ;
 PATH 372.4 357 372.4 381 ;
 END
END H PIN VDD DIRECTION INOUT ;
 SHAPE RING ;
 PORT LAYER M1 ;
 WIDTH 3.6 ;
 PATH 668 3.5 668 80.5 ;
 PATH 467 80.5 467 465.5 ;
 PATH 668 465.5 668 500.5 ;
 PATH 4 500.5 4 465.5 ;
 PATH 138 465.5 138 80.5 ;
 PATH 4 80.5 4 3.5 ;
 LAYER M2 ;
 WIDTH 3.6 ;
 PATH 4 3.5 668 3.5;
 PATH 668 80.5 467 80.5 ;
 PATH 467 465.5 668 465.5 ;
 PATH 668 500.5 4 500.5 ;
 PATH 4 465.5 138 465.5 ;
 PATH 138 80.5 4 80.5 ;
 END
END VDD PIN VSS DIRECTION INOUT ;
 SHAPE RING ;
 PORT LAYER M1 ;
 WIDTH 3.6 ;
 PATH 662 10 662 74 ;
 PATH 461 74 461 472 ;
 PATH 662 472 662 494 ;
 PATH 10 494 10 472;
 PATH 144 472 144 74 ;
 PATH 10 74 10 10 ;
LAYER M2 ;
 WIDTH 3.6 ;
 PATH 10 10 662 10 ;
 PATH 662 74 461 74 ;
 PATH 461 472 662 472 ;
 PATH 662 494 10 494 ;
 PATH 10 472 144 472 ;
 PATH 144 74 10 74 ;
 END
END VSS OBS LAYER M1 ;
 RECT 14 14 658 70 ;
 RECT 14 476 658 490 ;
 RECT 148 14 457 490 ;
 # rectilinear shape description LAYER OVERLAP ;
 RECT 0 0 672 84 ;
 RECT 134.4 84 470.4 462 ;
 RECT 0 462 672 504 ;
 END
END I2BLOCK 
