VIARULE VIALIST23
 LAYER M3 ;
 DIRECTION VERTICAL ;
 WIDTH 3.6 TO 3.6 ;
 LAYER M2 ;
 DIRECTION HORIZONTAL ;
 WIDTH 3.0 TO 3.0 ;
 VIA VIACENTER23 ;
 VIA VIATOP23 ;
 VIA VIABOTTOM23 ;
 VIA VIALEFT23 ;
 VIA VIARIGHT23 ;
END VIALIST23 
