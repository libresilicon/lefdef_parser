VIA C2NW DEFAULT
 LAYER NW ;
 RECT -2.0 -2.0 2.0 2.0 ;
 LAYER CUT01 ;
 RECT -0.6 -0.6 0.6 0.6 ;
 LAYER M1 ;
 RECT -2.0 -2.0 2.0 2.0 ;
END C2NW
